
module poly(I1,I2,I3,I4,I5,I6,O1);
  input  [11:0] I1;
  input  [11:0] I2;
  input  [11:0] I3;
  input [21:0] I4;
  input [21:0] I5;
  input [21:0] I6;

  output O1;

  wire [23:0] var_16 = {2'b00,I4};
  wire [23:0] var_17 = {2'b00,I5};
  wire [23:0] var_18 = {2'b00,I6};
  wire [13:0] var_12 = {2'b00,I1};
  wire [13:0] var_13 = {2'b00,I2};
  wire [13:0] var_14 = {2'b00,I3};
  wire [28:0] var_10 = {27'b000000000000000000000000000,2'b01};
  wire [23:0] var_19 = ((var_16 + var_17) + var_18);
  wire [27:0] var_15 = {14'b00000000000000,((var_12 + var_13) + var_14)};
  wire [28:0] var_11 = {15'b000000000000000,((14'b00000000000001 * var_14) + ((14'b00000000000001 * var_13) + ((14'b00000000000001 * var_12) + 14'b00000000000000)))};
  wire [26:0] tmp_0 = {3'b000,((24'b000000000000000000000001 * var_18) + ((24'b000000000000000000000001 * var_17) + ((24'b000000000000000000000001 * var_16) + 24'b000000000000000000000000)))};
  wire [26:0] tmp_1 = {25'b0000000000000000000000000,2'b11};
  wire tmp_2 = (tmp_0 < tmp_1);
  wire [28:0] tmp_3 = (((-{2'b00,tmp_2}) * var_10) + (((-{7'b0000000,I4}) * var_10) + (((-{7'b0000000,I5}) * var_10) + (((-{7'b0000000,I6}) * var_10) + ((var_11 * var_11) + 29'b00000000000000000000000000000)))));
  wire [27:0] tmp_4 = (var_15 * var_15);
  wire [27:0] tmp_5 = ({{{{1'b0,var_19},1'b0},1'b0},1'b0} + {{{{1'b0,1'b0},1'b0},1'b0},var_19});
  wire tmp_6 = (tmp_4 < tmp_5);
  wire lhs1 = ((tmp_3[28:28]) == (1'b1));
  wire rhs1 = tmp_6;

  assign O1 = (lhs1 == rhs1);

endmodule
