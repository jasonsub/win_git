
module mipsE ( clk, reset, memdata, memread, memwrite, adr, writedata, VMemr, 
        SMeml, VMeml, SMemr );
  input [7:0] memdata;
  output [7:0] adr;
  output [7:0] writedata;
  input clk, reset, VMemr, SMeml;
  output memread, memwrite, VMeml, SMemr;
  wire   pcen, VI1, alucont_2_, cont_SCI1, cont_VCint, cont_state_0_,
         cont_state_1_, cont_state_2_, cont_state_3_, dp_SABCI4P2, dp_VL,
         dp_aluout_0_, dp_aluout_1_, dp_aluout_2_, dp_aluout_3_, dp_aluout_4_,
         dp_aluout_5_, dp_aluout_6_, dp_aluout_7_, dp_aluresult_0_,
         dp_aluresult_1_, dp_aluresult_2_, dp_aluresult_3_, dp_aluresult_4_,
         dp_aluresult_5_, dp_aluresult_6_, dp_aluresult_7_, dp_SCI2I3LM2,
         dp_VB, dp_SCI2I3LM1, dp_VA, dp_SX2, dp_VM, dp_SABCI4LP, dp_VP,
         dp_pc_0_, dp_pc_1_, dp_pc_2_, dp_pc_3_, dp_pc_4_, dp_pc_5_, dp_pc_6_,
         dp_pc_7_, dp_SCX1, dp_SCX2, dp_VI2, dp_SCX3, dp_VI3, dp_SCX4, dp_VI4,
         cont_FCint_c, cont_FCint_e, cont_FCint_d, dp_rfE_RAM_0__0_,
         dp_rfE_RAM_0__1_, dp_rfE_RAM_0__2_, dp_rfE_RAM_0__3_,
         dp_rfE_RAM_0__4_, dp_rfE_RAM_0__5_, dp_rfE_RAM_0__6_,
         dp_rfE_RAM_0__7_, dp_rfE_RAM_1__0_, dp_rfE_RAM_1__1_,
         dp_rfE_RAM_1__2_, dp_rfE_RAM_1__3_, dp_rfE_RAM_1__4_,
         dp_rfE_RAM_1__5_, dp_rfE_RAM_1__6_, dp_rfE_RAM_1__7_,
         dp_rfE_RAM_2__0_, dp_rfE_RAM_2__1_, dp_rfE_RAM_2__2_,
         dp_rfE_RAM_2__3_, dp_rfE_RAM_2__4_, dp_rfE_RAM_2__5_,
         dp_rfE_RAM_2__6_, dp_rfE_RAM_2__7_, dp_rfE_RAM_3__0_,
         dp_rfE_RAM_3__1_, dp_rfE_RAM_3__2_, dp_rfE_RAM_3__3_,
         dp_rfE_RAM_3__4_, dp_rfE_RAM_3__5_, dp_rfE_RAM_3__6_,
         dp_rfE_RAM_3__7_, dp_rfE_RAM_4__0_, dp_rfE_RAM_4__1_,
         dp_rfE_RAM_4__2_, dp_rfE_RAM_4__3_, dp_rfE_RAM_4__4_,
         dp_rfE_RAM_4__5_, dp_rfE_RAM_4__6_, dp_rfE_RAM_4__7_,
         dp_rfE_RAM_5__0_, dp_rfE_RAM_5__1_, dp_rfE_RAM_5__2_,
         dp_rfE_RAM_5__3_, dp_rfE_RAM_5__4_, dp_rfE_RAM_5__5_,
         dp_rfE_RAM_5__6_, dp_rfE_RAM_5__7_, dp_rfE_RAM_6__0_,
         dp_rfE_RAM_6__1_, dp_rfE_RAM_6__2_, dp_rfE_RAM_6__3_,
         dp_rfE_RAM_6__4_, dp_rfE_RAM_6__5_, dp_rfE_RAM_6__6_,
         dp_rfE_RAM_6__7_, dp_rfE_RAM_7__0_, dp_rfE_RAM_7__1_,
         dp_rfE_RAM_7__2_, dp_rfE_RAM_7__3_, dp_rfE_RAM_7__4_,
         dp_rfE_RAM_7__5_, dp_rfE_RAM_7__6_, dp_rfE_RAM_7__7_,
         dp_alunit_sum_0_, dp_alunit_sum_1_, dp_alunit_sum_2_,
         dp_alunit_sum_3_, dp_alunit_sum_4_, dp_alunit_sum_5_,
         dp_alunit_sum_6_, dp_alunit_sum_7_, dp_FB_c, dp_FB_b, dp_FB_e,
         dp_FB_d, dp_FP_c, dp_FP_e, dp_FP_d, dp_FCI2I3LM_c, dp_FCI2I3LM_b,
         dp_FCI2I3LM_e, dp_FCI2I3LM_d, dp_FABCI4P_c, dp_FABCI4P_b,
         dp_FABCI4P_e, dp_FX_c, dp_FX_b, dp_FX_e, dp_FX_d, dp_EBREnP_Es,
         cont_EBRC_eBCtl1_d, cont_EBRC_eBCtl1_e, cont_EBRC_eBCtl1_b,
         cont_EBRC_eBCtl1_f, cont_FCint_pDFFS1_qi, dp_FL_EFork22_c,
         dp_FL_EFork22_e, dp_FL_EFork22_d, dp_FL_EFork21_c, dp_FL_EFork21_b,
         dp_FL_EFork21_e, dp_FCX_EFork21_c, dp_FCX_EFork21_b, dp_FCX_EFork21_e,
         dp_FCX_EFork21_d, dp_FC_EFork21_c, dp_FC_EFork21_b, dp_FC_EFork21_e,
         dp_FC_EFork21_d, dp_EBL_eBCtl1_d, dp_EBL_eBCtl1_e, dp_EBL_eBCtl1_b,
         dp_EBL_eBCtl1_f, dp_EBB_eBCtl1_d, dp_EBB_eBCtl1_e, dp_EBB_eBCtl1_b,
         dp_EBB_eBCtl1_f, dp_EBA_eBCtl1_d, dp_EBA_eBCtl1_e, dp_EBA_eBCtl1_b,
         dp_EBA_eBCtl1_f, dp_EBM_eBCtl1_d, dp_EBM_eBCtl1_e, dp_EBM_eBCtl1_b,
         dp_EBM_eBCtl1_f, dp_EBREnP_eBCtl1_d, dp_EBREnP_eBCtl1_e,
         dp_EBREnP_eBCtl1_b, dp_EBREnP_eBCtl1_f, dp_EBREnI1_eBCtl1_d,
         dp_EBREnI1_eBCtl1_e, dp_EBREnI1_eBCtl1_b, dp_EBREnI1_eBCtl1_f,
         dp_EBREnI2_eBCtl1_d, dp_EBREnI2_eBCtl1_e, dp_EBREnI2_eBCtl1_b,
         dp_EBREnI2_eBCtl1_f, dp_EBREnI3_eBCtl1_d, dp_EBREnI3_eBCtl1_e,
         dp_EBREnI3_eBCtl1_b, dp_EBREnI3_eBCtl1_f, dp_EBREnI4_eBCtl1_d,
         dp_EBREnI4_eBCtl1_e, dp_EBREnI4_eBCtl1_b, dp_EBREnI4_eBCtl1_f,
         dp_FB_pDFFS0_qi, dp_FB_pDFFS1_qi, dp_FP_pDFFS0_qi, dp_FP_pDFFS1_qi,
         dp_FCI2I3LM_pDFFS0_qi, dp_FCI2I3LM_pDFFS1_qi, dp_FABCI4P_pDFFS0_qi,
         dp_FABCI4P_pDFFS1_qi, dp_FX_pDFFS0_qi, dp_FX_pDFFS1_qi,
         cont_FCint_pDFFS0_qi, cont_EBRC_eBCtl1_iLHS1_di,
         cont_EBRC_eBCtl1_iLLS2_di, dp_FCX_EFork31_EFork22_c,
         dp_FCX_EFork31_EFork22_b, dp_FCX_EFork31_EFork22_e,
         dp_FCX_EFork31_EFork22_d, dp_FCX_EFork31_EFork21_c,
         dp_FCX_EFork31_EFork21_b, dp_FCX_EFork31_EFork21_e,
         dp_FCX_EFork31_EFork21_d, dp_FC_EFork31_EFork22_c,
         dp_FC_EFork31_EFork22_b, dp_FC_EFork31_EFork22_e,
         dp_FC_EFork31_EFork22_d, dp_FC_EFork31_EFork21_c,
         dp_FC_EFork31_EFork21_e, dp_FC_EFork31_EFork21_d,
         dp_FL_EFork22_pDFFS0_qi, dp_FL_EFork22_pDFFS1_qi,
         dp_FL_EFork21_pDFFS0_qi, dp_FL_EFork21_pDFFS1_qi,
         dp_FCX_EFork21_pDFFS0_qi, dp_FCX_EFork21_pDFFS1_qi,
         dp_FC_EFork21_pDFFS0_qi, dp_FC_EFork21_pDFFS1_qi,
         cont_EBRC_lLRE1_U3_clki, cont_EBRC_lHRE1_U3_clki, dp_FB_pDFFS0_U1_di,
         dp_FB_pDFFS1_U1_di, dp_FP_pDFFS0_U1_di, dp_FP_pDFFS1_U1_di,
         dp_FCI2I3LM_pDFFS0_U1_di, dp_FCI2I3LM_pDFFS1_U1_di,
         dp_FABCI4P_pDFFS0_U1_di, dp_FABCI4P_pDFFS1_U1_di, dp_FX_pDFFS0_U1_di,
         dp_FX_pDFFS1_U1_di, dp_EBL_eBCtl1_iLHS1_di, dp_EBB_eBCtl1_iLHS1_di,
         dp_EBA_eBCtl1_iLHS1_di, dp_EBM_eBCtl1_iLHS1_di,
         dp_EBREnP_eBCtl1_iLHS1_di, dp_EBREnI1_eBCtl1_iLHS1_di,
         dp_EBREnI2_eBCtl1_iLHS1_di, dp_EBREnI3_eBCtl1_iLHS1_di,
         dp_EBREnI4_eBCtl1_iLHS1_di, cont_FCint_pDFFS0_U1_di,
         cont_FCint_pDFFS1_U1_di, dp_EBL_eBCtl1_iLLS2_di,
         dp_EBB_eBCtl1_iLLS2_di, dp_EBA_eBCtl1_iLLS2_di,
         dp_EBM_eBCtl1_iLLS2_di, dp_EBREnP_eBCtl1_iLLS2_di,
         dp_EBREnI1_eBCtl1_iLLS2_di, dp_EBREnI2_eBCtl1_iLLS2_di,
         dp_EBREnI3_eBCtl1_iLLS2_di, dp_EBREnI4_eBCtl1_iLLS2_di,
         dp_EBREnP_U0_U7_clki, dp_EBREnI1_U0_U7_clki, dp_EBREnI2_U0_U7_clki,
         dp_EBREnI3_U0_U5_clki, dp_EBREnI4_U0_U7_clki, dp_EBREnP_U1_U7_clki,
         dp_EBREnP_U1_U6_clki, dp_EBREnP_U1_U5_clki, dp_EBREnP_U1_U4_clki,
         dp_EBREnP_U1_U3_clki, dp_EBREnP_U1_U2_clki, dp_EBREnP_U1_U1_clki,
         dp_EBREnP_U1_U0_clki, dp_EBREnI1_U1_U7_clki, dp_EBREnI2_U1_U7_clki,
         dp_EBREnI3_U1_U5_clki, dp_EBREnI4_U1_U7_clki, dp_EBL_U0_U7_clki,
         dp_EBB_U0_U7_clki, dp_EBA_U0_U7_clki, dp_EBM_U0_U7_clki,
         dp_EBL_U1_U7_clki, dp_EBB_U1_U7_clki, dp_EBA_U1_U7_clki,
         dp_EBM_U1_U7_clki, dp_FCX_EFork31_EFork22_pDFFS0_qi,
         dp_FCX_EFork31_EFork22_pDFFS1_qi, dp_FCX_EFork31_EFork21_pDFFS0_qi,
         dp_FCX_EFork31_EFork21_pDFFS1_qi, dp_FC_EFork31_EFork22_pDFFS0_qi,
         dp_FC_EFork31_EFork22_pDFFS1_qi, dp_FC_EFork31_EFork21_pDFFS0_qi,
         dp_FC_EFork31_EFork21_pDFFS1_qi, dp_FL_EFork22_pDFFS0_U1_di,
         dp_FL_EFork22_pDFFS1_U1_di, dp_FL_EFork21_pDFFS0_U1_di,
         dp_FL_EFork21_pDFFS1_U1_di, dp_FCX_EFork21_pDFFS0_U1_di,
         dp_FCX_EFork21_pDFFS1_U1_di, dp_FC_EFork21_pDFFS0_U1_di,
         dp_FC_EFork21_pDFFS1_U1_di, dp_FCX_EFork31_EFork22_pDFFS0_U1_di,
         dp_FCX_EFork31_EFork22_pDFFS1_U1_di,
         dp_FCX_EFork31_EFork21_pDFFS0_U1_di,
         dp_FCX_EFork31_EFork21_pDFFS1_U1_di,
         dp_FC_EFork31_EFork22_pDFFS0_U1_di,
         dp_FC_EFork31_EFork22_pDFFS1_U1_di,
         dp_FC_EFork31_EFork21_pDFFS0_U1_di,
         dp_FC_EFork31_EFork21_pDFFS1_U1_di, n65, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n94, n95, n96, n97, n98, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n1, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, DP_OP_50_64_8725_n85,
         DP_OP_50_64_8725_n71, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753;
  wire   [31:0] instr;
  wire   [3:0] cont_nextstate;
  wire   [7:0] dp_src1;
  wire   [7:0] dp_rd2;
  wire   [7:0] dp_a;
  wire   [7:0] dp_rd1;
  wire   [7:0] dp_md;
  wire   [7:0] dp_nextpc;
  wire   [3:0] cont_EBRC_m;
  wire   [7:0] dp_EBREnI4_m;
  wire   [7:0] dp_EBM_m;
  wire   [7:0] dp_alunit_b2;
  wire   [7:0] dp_EBREnP_m;
  wire   [7:0] dp_EBREnI1_m;
  wire   [7:0] dp_EBREnI2_m;
  wire   [7:0] dp_EBREnI3_m;
  wire   [7:0] dp_EBL_m;
  wire   [7:0] dp_EBB_m;
  wire   [7:0] dp_EBA_m;

  LCX1 cont_EBRC_lLRE1_U0_U4 ( .CLR(n753), .G(cont_EBRC_lLRE1_U3_clki), .D(
        cont_nextstate[0]), .Q(cont_EBRC_m[0]) );
  LCNX1 cont_EBRC_lHRE1_U0_U3 ( .CLR(n752), .D(cont_EBRC_m[0]), .G(
        cont_EBRC_lHRE1_U3_clki), .Q(cont_state_0_) );
  LCX1 cont_EBRC_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(
        cont_EBRC_eBCtl1_iLHS1_di), .Q(cont_VCint) );
  LCX1 cont_EBRC_eBCtl1_iLHR1_U1 ( .CLR(n753), .G(clk), .D(cont_EBRC_eBCtl1_f), 
        .Q(cont_SCI1) );
  LCNX1 cont_EBRC_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(cont_EBRC_eBCtl1_iLLS2_di), 
        .G(clk), .Q(cont_EBRC_eBCtl1_b) );
  LCNX1 cont_EBRC_eBCtl1_iLLR2_U1 ( .CLR(n752), .D(cont_EBRC_eBCtl1_e), .G(clk), .Q(cont_EBRC_eBCtl1_d) );
  LCX1 dp_EBREnI4_U0_U0_U4 ( .CLR(n753), .G(dp_EBREnI4_U0_U7_clki), .D(
        memdata[0]), .Q(dp_EBREnI4_m[0]) );
  LCNX1 dp_EBREnI4_U1_U0_U3 ( .CLR(n752), .D(dp_EBREnI4_m[0]), .G(
        dp_EBREnI4_U1_U7_clki), .Q(instr[0]) );
  LCX1 dp_EBM_U0_U0_U4 ( .CLR(n1), .G(dp_EBM_U0_U7_clki), .D(memdata[0]), .Q(
        dp_EBM_m[0]) );
  LCNX1 dp_EBM_U1_U0_U3 ( .CLR(n1), .D(dp_EBM_m[0]), .G(dp_EBM_U1_U7_clki), 
        .Q(dp_md[0]) );
  LCX1 cont_EBRC_lLRE1_U3_U4 ( .CLR(n753), .G(cont_EBRC_lLRE1_U3_clki), .D(
        cont_nextstate[3]), .Q(cont_EBRC_m[3]) );
  LCX1 cont_EBRC_lLRE1_U2_U4 ( .CLR(n753), .G(cont_EBRC_lLRE1_U3_clki), .D(
        cont_nextstate[2]), .Q(cont_EBRC_m[2]) );
  LCX1 cont_EBRC_lLRE1_U1_U4 ( .CLR(n753), .G(cont_EBRC_lLRE1_U3_clki), .D(
        cont_nextstate[1]), .Q(cont_EBRC_m[1]) );
  LCNX1 cont_EBRC_lHRE1_U3_U3 ( .CLR(n752), .D(cont_EBRC_m[3]), .G(
        cont_EBRC_lHRE1_U3_clki), .Q(cont_state_3_) );
  LCNX1 cont_EBRC_lHRE1_U2_U3 ( .CLR(n752), .D(cont_EBRC_m[2]), .G(
        cont_EBRC_lHRE1_U3_clki), .Q(cont_state_2_) );
  LCNX1 cont_EBRC_lHRE1_U1_U3 ( .CLR(n752), .D(cont_EBRC_m[1]), .G(
        cont_EBRC_lHRE1_U3_clki), .Q(cont_state_1_) );
  LCX1 dp_FB_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(dp_FB_pDFFS0_U1_di), .Q(
        dp_FB_c) );
  LCX1 dp_FB_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(dp_FB_pDFFS1_U1_di), .Q(
        dp_FB_e) );
  LCX1 dp_FP_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(dp_FP_pDFFS0_U1_di), .Q(
        dp_FP_c) );
  LCX1 dp_FP_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(dp_FP_pDFFS1_U1_di), .Q(
        dp_FP_e) );
  LCX1 dp_FCI2I3LM_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FCI2I3LM_pDFFS0_U1_di), .Q(dp_FCI2I3LM_c) );
  LCX1 dp_FCI2I3LM_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FCI2I3LM_pDFFS1_U1_di), .Q(dp_FCI2I3LM_e) );
  LCX1 dp_FABCI4P_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(dp_FABCI4P_pDFFS0_U1_di), .Q(dp_FABCI4P_c) );
  LCX1 dp_FABCI4P_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(dp_FABCI4P_pDFFS1_U1_di), .Q(dp_FABCI4P_e) );
  LCX1 dp_FX_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(dp_FX_pDFFS0_U1_di), .Q(
        dp_FX_c) );
  LCX1 dp_FX_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(dp_FX_pDFFS1_U1_di), .Q(
        dp_FX_e) );
  LCX1 dp_EBL_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(dp_EBL_eBCtl1_iLHS1_di), 
        .Q(dp_VL) );
  LCX1 dp_EBB_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(dp_EBB_eBCtl1_iLHS1_di), 
        .Q(dp_VB) );
  LCX1 dp_EBA_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(dp_EBA_eBCtl1_iLHS1_di), 
        .Q(dp_VA) );
  LCX1 dp_EBM_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(dp_EBM_eBCtl1_iLHS1_di), 
        .Q(dp_VM) );
  LCX1 dp_EBREnP_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(
        dp_EBREnP_eBCtl1_iLHS1_di), .Q(dp_VP) );
  LCX1 dp_EBREnI1_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(
        dp_EBREnI1_eBCtl1_iLHS1_di), .Q(VI1) );
  LCX1 dp_EBREnI2_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(
        dp_EBREnI2_eBCtl1_iLHS1_di), .Q(dp_VI2) );
  LCX1 dp_EBREnI3_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(
        dp_EBREnI3_eBCtl1_iLHS1_di), .Q(dp_VI3) );
  LCX1 dp_EBREnI4_eBCtl1_iLHS1_U3 ( .CLR(n1), .G(clk), .D(
        dp_EBREnI4_eBCtl1_iLHS1_di), .Q(dp_VI4) );
  LCX1 cont_FCint_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(cont_FCint_pDFFS0_U1_di), .Q(cont_FCint_c) );
  LCX1 cont_FCint_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(cont_FCint_pDFFS1_U1_di), .Q(cont_FCint_e) );
  LCX1 dp_EBL_eBCtl1_iLHR1_U1 ( .CLR(n581), .G(clk), .D(dp_EBL_eBCtl1_f), .Q(
        dp_SABCI4P2) );
  LCX1 dp_EBB_eBCtl1_iLHR1_U1 ( .CLR(n753), .G(clk), .D(dp_EBB_eBCtl1_f), .Q(
        dp_SCI2I3LM2) );
  LCX1 dp_EBA_eBCtl1_iLHR1_U1 ( .CLR(n581), .G(clk), .D(dp_EBA_eBCtl1_f), .Q(
        dp_SCI2I3LM1) );
  LCX1 dp_EBM_eBCtl1_iLHR1_U1 ( .CLR(n581), .G(clk), .D(dp_EBM_eBCtl1_f), .Q(
        dp_SX2) );
  LCX1 dp_EBREnP_eBCtl1_iLHR1_U1 ( .CLR(n581), .G(clk), .D(dp_EBREnP_eBCtl1_f), 
        .Q(dp_SABCI4LP) );
  LCX1 dp_EBREnI1_eBCtl1_iLHR1_U1 ( .CLR(n581), .G(clk), .D(
        dp_EBREnI1_eBCtl1_f), .Q(dp_SCX1) );
  LCX1 dp_EBREnI2_eBCtl1_iLHR1_U1 ( .CLR(n581), .G(clk), .D(
        dp_EBREnI2_eBCtl1_f), .Q(dp_SCX2) );
  LCX1 dp_EBREnI3_eBCtl1_iLHR1_U1 ( .CLR(n581), .G(clk), .D(
        dp_EBREnI3_eBCtl1_f), .Q(dp_SCX3) );
  LCX1 dp_EBREnI4_eBCtl1_iLHR1_U1 ( .CLR(n581), .G(clk), .D(
        dp_EBREnI4_eBCtl1_f), .Q(dp_SCX4) );
  LCNX1 dp_EBL_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBL_eBCtl1_iLLS2_di), .G(clk), 
        .Q(dp_EBL_eBCtl1_b) );
  LCNX1 dp_EBB_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBB_eBCtl1_iLLS2_di), .G(clk), 
        .Q(dp_EBB_eBCtl1_b) );
  LCNX1 dp_EBA_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBA_eBCtl1_iLLS2_di), .G(clk), 
        .Q(dp_EBA_eBCtl1_b) );
  LCNX1 dp_EBM_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBM_eBCtl1_iLLS2_di), .G(clk), 
        .Q(dp_EBM_eBCtl1_b) );
  LCNX1 dp_EBREnP_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBREnP_eBCtl1_iLLS2_di), 
        .G(clk), .Q(dp_EBREnP_eBCtl1_b) );
  LCNX1 dp_EBREnI1_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBREnI1_eBCtl1_iLLS2_di), 
        .G(clk), .Q(dp_EBREnI1_eBCtl1_b) );
  LCNX1 dp_EBREnI2_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBREnI2_eBCtl1_iLLS2_di), 
        .G(clk), .Q(dp_EBREnI2_eBCtl1_b) );
  LCNX1 dp_EBREnI3_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBREnI3_eBCtl1_iLLS2_di), 
        .G(clk), .Q(dp_EBREnI3_eBCtl1_b) );
  LCNX1 dp_EBREnI4_eBCtl1_iLLS2_U3 ( .CLR(n1), .D(dp_EBREnI4_eBCtl1_iLLS2_di), 
        .G(clk), .Q(dp_EBREnI4_eBCtl1_b) );
  LCNX1 dp_FB_pDFFS0_U0_U1 ( .CLR(n752), .D(dp_FB_b), .G(clk), .Q(
        dp_FB_pDFFS0_qi) );
  LCNX1 dp_FB_pDFFS1_U0_U1 ( .CLR(n752), .D(dp_FB_d), .G(clk), .Q(
        dp_FB_pDFFS1_qi) );
  LCNX1 dp_FP_pDFFS0_U0_U1 ( .CLR(n752), .D(n75), .G(clk), .Q(dp_FP_pDFFS0_qi)
         );
  LCNX1 dp_FP_pDFFS1_U0_U1 ( .CLR(n753), .D(dp_FP_d), .G(clk), .Q(
        dp_FP_pDFFS1_qi) );
  LCNX1 dp_FCI2I3LM_pDFFS0_U0_U1 ( .CLR(n753), .D(dp_FCI2I3LM_b), .G(clk), .Q(
        dp_FCI2I3LM_pDFFS0_qi) );
  LCNX1 dp_FCI2I3LM_pDFFS1_U0_U1 ( .CLR(n753), .D(dp_FCI2I3LM_d), .G(clk), .Q(
        dp_FCI2I3LM_pDFFS1_qi) );
  LCNX1 dp_FABCI4P_pDFFS0_U0_U1 ( .CLR(n753), .D(dp_FABCI4P_b), .G(clk), .Q(
        dp_FABCI4P_pDFFS0_qi) );
  LCNX1 dp_FABCI4P_pDFFS1_U0_U1 ( .CLR(n753), .D(n130), .G(clk), .Q(
        dp_FABCI4P_pDFFS1_qi) );
  LCNX1 dp_FX_pDFFS0_U0_U1 ( .CLR(n753), .D(dp_FX_b), .G(clk), .Q(
        dp_FX_pDFFS0_qi) );
  LCNX1 dp_FX_pDFFS1_U0_U1 ( .CLR(n753), .D(dp_FX_d), .G(clk), .Q(
        dp_FX_pDFFS1_qi) );
  LCNX1 dp_EBL_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBL_eBCtl1_e), .G(clk), .Q(
        dp_EBL_eBCtl1_d) );
  LCNX1 dp_EBB_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBB_eBCtl1_e), .G(clk), .Q(
        dp_EBB_eBCtl1_d) );
  LCNX1 dp_EBA_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBA_eBCtl1_e), .G(clk), .Q(
        dp_EBA_eBCtl1_d) );
  LCNX1 dp_EBM_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBM_eBCtl1_e), .G(clk), .Q(
        dp_EBM_eBCtl1_d) );
  LCNX1 dp_EBREnP_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBREnP_eBCtl1_e), .G(clk), .Q(dp_EBREnP_eBCtl1_d) );
  LCNX1 dp_EBREnI1_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBREnI1_eBCtl1_e), .G(
        clk), .Q(dp_EBREnI1_eBCtl1_d) );
  LCNX1 dp_EBREnI2_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBREnI2_eBCtl1_e), .G(
        clk), .Q(dp_EBREnI2_eBCtl1_d) );
  LCNX1 dp_EBREnI3_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBREnI3_eBCtl1_e), .G(
        clk), .Q(dp_EBREnI3_eBCtl1_d) );
  LCNX1 dp_EBREnI4_eBCtl1_iLLR2_U1 ( .CLR(n753), .D(dp_EBREnI4_eBCtl1_e), .G(
        clk), .Q(dp_EBREnI4_eBCtl1_d) );
  LCNX1 cont_FCint_pDFFS0_U0_U1 ( .CLR(n753), .D(n69), .G(clk), .Q(
        cont_FCint_pDFFS0_qi) );
  LCNX1 cont_FCint_pDFFS1_U0_U1 ( .CLR(n753), .D(cont_FCint_d), .G(clk), .Q(
        cont_FCint_pDFFS1_qi) );
  LCX1 dp_EBREnP_U0_U7_U4 ( .CLR(n581), .G(dp_EBREnP_U0_U7_clki), .D(
        dp_nextpc[7]), .Q(dp_EBREnP_m[7]) );
  LCX1 dp_EBREnP_U0_U6_U4 ( .CLR(n581), .G(dp_EBREnP_U0_U7_clki), .D(
        dp_nextpc[6]), .Q(dp_EBREnP_m[6]) );
  LCX1 dp_EBREnP_U0_U5_U4 ( .CLR(n753), .G(dp_EBREnP_U0_U7_clki), .D(
        dp_nextpc[5]), .Q(dp_EBREnP_m[5]) );
  LCX1 dp_EBREnP_U0_U4_U4 ( .CLR(n581), .G(dp_EBREnP_U0_U7_clki), .D(
        dp_nextpc[4]), .Q(dp_EBREnP_m[4]) );
  LCX1 dp_EBREnP_U0_U3_U4 ( .CLR(n581), .G(dp_EBREnP_U0_U7_clki), .D(
        dp_nextpc[3]), .Q(dp_EBREnP_m[3]) );
  LCX1 dp_EBREnP_U0_U2_U4 ( .CLR(n581), .G(dp_EBREnP_U0_U7_clki), .D(
        dp_nextpc[2]), .Q(dp_EBREnP_m[2]) );
  LCX1 dp_EBREnP_U0_U1_U4 ( .CLR(n581), .G(dp_EBREnP_U0_U7_clki), .D(n100), 
        .Q(dp_EBREnP_m[1]) );
  LCX1 dp_EBREnP_U0_U0_U4 ( .CLR(n581), .G(dp_EBREnP_U0_U7_clki), .D(n98), .Q(
        dp_EBREnP_m[0]) );
  LCX1 dp_EBREnI1_U0_U7_U4 ( .CLR(n581), .G(dp_EBREnI1_U0_U7_clki), .D(
        memdata[7]), .Q(dp_EBREnI1_m[7]) );
  LCX1 dp_EBREnI1_U0_U6_U4 ( .CLR(n581), .G(dp_EBREnI1_U0_U7_clki), .D(
        memdata[6]), .Q(dp_EBREnI1_m[6]) );
  LCX1 dp_EBREnI1_U0_U5_U4 ( .CLR(n581), .G(dp_EBREnI1_U0_U7_clki), .D(
        memdata[5]), .Q(dp_EBREnI1_m[5]) );
  LCX1 dp_EBREnI1_U0_U4_U4 ( .CLR(n581), .G(dp_EBREnI1_U0_U7_clki), .D(
        memdata[4]), .Q(dp_EBREnI1_m[4]) );
  LCX1 dp_EBREnI1_U0_U3_U4 ( .CLR(n581), .G(dp_EBREnI1_U0_U7_clki), .D(
        memdata[3]), .Q(dp_EBREnI1_m[3]) );
  LCX1 dp_EBREnI1_U0_U2_U4 ( .CLR(n581), .G(dp_EBREnI1_U0_U7_clki), .D(
        memdata[2]), .Q(dp_EBREnI1_m[2]) );
  LCX1 dp_EBREnI2_U0_U7_U4 ( .CLR(n581), .G(dp_EBREnI2_U0_U7_clki), .D(
        memdata[7]), .Q(dp_EBREnI2_m[7]) );
  LCX1 dp_EBREnI2_U0_U6_U4 ( .CLR(n581), .G(dp_EBREnI2_U0_U7_clki), .D(
        memdata[6]), .Q(dp_EBREnI2_m[6]) );
  LCX1 dp_EBREnI2_U0_U5_U4 ( .CLR(n581), .G(dp_EBREnI2_U0_U7_clki), .D(
        memdata[5]), .Q(dp_EBREnI2_m[5]) );
  LCX1 dp_EBREnI2_U0_U2_U4 ( .CLR(n581), .G(dp_EBREnI2_U0_U7_clki), .D(
        memdata[2]), .Q(dp_EBREnI2_m[2]) );
  LCX1 dp_EBREnI2_U0_U1_U4 ( .CLR(n581), .G(dp_EBREnI2_U0_U7_clki), .D(
        memdata[1]), .Q(dp_EBREnI2_m[1]) );
  LCX1 dp_EBREnI2_U0_U0_U4 ( .CLR(n581), .G(dp_EBREnI2_U0_U7_clki), .D(
        memdata[0]), .Q(dp_EBREnI2_m[0]) );
  LCX1 dp_EBREnI3_U0_U5_U4 ( .CLR(n581), .G(dp_EBREnI3_U0_U5_clki), .D(
        memdata[5]), .Q(dp_EBREnI3_m[5]) );
  LCX1 dp_EBREnI3_U0_U4_U4 ( .CLR(n581), .G(dp_EBREnI3_U0_U5_clki), .D(
        memdata[4]), .Q(dp_EBREnI3_m[4]) );
  LCX1 dp_EBREnI3_U0_U3_U4 ( .CLR(n581), .G(dp_EBREnI3_U0_U5_clki), .D(
        memdata[3]), .Q(dp_EBREnI3_m[3]) );
  LCX1 dp_EBREnI4_U0_U7_U4 ( .CLR(n581), .G(dp_EBREnI4_U0_U7_clki), .D(
        memdata[7]), .Q(dp_EBREnI4_m[7]) );
  LCX1 dp_EBREnI4_U0_U6_U4 ( .CLR(n581), .G(dp_EBREnI4_U0_U7_clki), .D(
        memdata[6]), .Q(dp_EBREnI4_m[6]) );
  LCX1 dp_EBREnI4_U0_U5_U4 ( .CLR(n581), .G(dp_EBREnI4_U0_U7_clki), .D(
        memdata[5]), .Q(dp_EBREnI4_m[5]) );
  LCX1 dp_EBREnI4_U0_U4_U4 ( .CLR(n581), .G(dp_EBREnI4_U0_U7_clki), .D(
        memdata[4]), .Q(dp_EBREnI4_m[4]) );
  LCX1 dp_EBREnI4_U0_U3_U4 ( .CLR(n581), .G(dp_EBREnI4_U0_U7_clki), .D(
        memdata[3]), .Q(dp_EBREnI4_m[3]) );
  LCX1 dp_EBREnI4_U0_U2_U4 ( .CLR(n581), .G(dp_EBREnI4_U0_U7_clki), .D(
        memdata[2]), .Q(dp_EBREnI4_m[2]) );
  LCX1 dp_EBREnI4_U0_U1_U4 ( .CLR(n753), .G(dp_EBREnI4_U0_U7_clki), .D(
        memdata[1]), .Q(dp_EBREnI4_m[1]) );
  LCNX1 dp_EBREnP_U1_U7_U3 ( .CLR(n753), .D(dp_EBREnP_m[7]), .G(
        dp_EBREnP_U1_U7_clki), .Q(dp_pc_7_) );
  NAND3X1 dp_EBREnP_U1_U7_U2 ( .A(pcen), .B(dp_EBREnP_Es), .C(clk), .Y(
        dp_EBREnP_U1_U7_clki) );
  LCNX1 dp_EBREnP_U1_U6_U3 ( .CLR(n753), .D(dp_EBREnP_m[6]), .G(
        dp_EBREnP_U1_U6_clki), .Q(dp_pc_6_) );
  NAND3X1 dp_EBREnP_U1_U6_U2 ( .A(pcen), .B(dp_EBREnP_Es), .C(clk), .Y(
        dp_EBREnP_U1_U6_clki) );
  LCNX1 dp_EBREnP_U1_U5_U3 ( .CLR(n753), .D(dp_EBREnP_m[5]), .G(
        dp_EBREnP_U1_U5_clki), .Q(dp_pc_5_) );
  NAND3X1 dp_EBREnP_U1_U5_U2 ( .A(pcen), .B(dp_EBREnP_Es), .C(clk), .Y(
        dp_EBREnP_U1_U5_clki) );
  LCNX1 dp_EBREnP_U1_U4_U3 ( .CLR(n753), .D(dp_EBREnP_m[4]), .G(
        dp_EBREnP_U1_U4_clki), .Q(dp_pc_4_) );
  NAND3X1 dp_EBREnP_U1_U4_U2 ( .A(pcen), .B(dp_EBREnP_Es), .C(clk), .Y(
        dp_EBREnP_U1_U4_clki) );
  LCNX1 dp_EBREnP_U1_U3_U3 ( .CLR(n753), .D(dp_EBREnP_m[3]), .G(
        dp_EBREnP_U1_U3_clki), .Q(dp_pc_3_) );
  NAND3X1 dp_EBREnP_U1_U3_U2 ( .A(pcen), .B(dp_EBREnP_Es), .C(clk), .Y(
        dp_EBREnP_U1_U3_clki) );
  LCNX1 dp_EBREnP_U1_U2_U3 ( .CLR(n753), .D(dp_EBREnP_m[2]), .G(
        dp_EBREnP_U1_U2_clki), .Q(dp_pc_2_) );
  NAND3X1 dp_EBREnP_U1_U2_U2 ( .A(pcen), .B(dp_EBREnP_Es), .C(clk), .Y(
        dp_EBREnP_U1_U2_clki) );
  LCNX1 dp_EBREnP_U1_U1_U3 ( .CLR(n753), .D(dp_EBREnP_m[1]), .G(
        dp_EBREnP_U1_U1_clki), .Q(dp_pc_1_) );
  NAND3X1 dp_EBREnP_U1_U1_U2 ( .A(pcen), .B(dp_EBREnP_Es), .C(clk), .Y(
        dp_EBREnP_U1_U1_clki) );
  LCNX1 dp_EBREnP_U1_U0_U3 ( .CLR(n753), .D(dp_EBREnP_m[0]), .G(
        dp_EBREnP_U1_U0_clki), .Q(dp_pc_0_) );
  NAND3X1 dp_EBREnP_U1_U0_U2 ( .A(pcen), .B(dp_EBREnP_Es), .C(clk), .Y(
        dp_EBREnP_U1_U0_clki) );
  LCNX1 dp_EBREnI1_U1_U7_U3 ( .CLR(n753), .D(dp_EBREnI1_m[7]), .G(
        dp_EBREnI1_U1_U7_clki), .Q(instr[31]) );
  LCNX1 dp_EBREnI1_U1_U6_U3 ( .CLR(n753), .D(dp_EBREnI1_m[6]), .G(
        dp_EBREnI1_U1_U7_clki), .Q(instr[30]) );
  LCNX1 dp_EBREnI1_U1_U5_U3 ( .CLR(n581), .D(dp_EBREnI1_m[5]), .G(
        dp_EBREnI1_U1_U7_clki), .Q(instr[29]) );
  LCNX1 dp_EBREnI1_U1_U4_U3 ( .CLR(n581), .D(dp_EBREnI1_m[4]), .G(
        dp_EBREnI1_U1_U7_clki), .Q(instr[28]) );
  LCNX1 dp_EBREnI1_U1_U3_U3 ( .CLR(n581), .D(dp_EBREnI1_m[3]), .G(
        dp_EBREnI1_U1_U7_clki), .Q(instr[27]) );
  LCNX1 dp_EBREnI1_U1_U2_U3 ( .CLR(n581), .D(dp_EBREnI1_m[2]), .G(
        dp_EBREnI1_U1_U7_clki), .Q(instr[26]) );
  LCNX1 dp_EBREnI2_U1_U7_U3 ( .CLR(n753), .D(dp_EBREnI2_m[7]), .G(
        dp_EBREnI2_U1_U7_clki), .Q(instr[23]) );
  LCNX1 dp_EBREnI2_U1_U6_U3 ( .CLR(n581), .D(dp_EBREnI2_m[6]), .G(
        dp_EBREnI2_U1_U7_clki), .Q(instr[22]) );
  LCNX1 dp_EBREnI2_U1_U5_U3 ( .CLR(n753), .D(dp_EBREnI2_m[5]), .G(
        dp_EBREnI2_U1_U7_clki), .Q(instr[21]) );
  LCNX1 dp_EBREnI2_U1_U2_U3 ( .CLR(n753), .D(dp_EBREnI2_m[2]), .G(
        dp_EBREnI2_U1_U7_clki), .Q(instr[18]) );
  LCNX1 dp_EBREnI2_U1_U1_U3 ( .CLR(n581), .D(dp_EBREnI2_m[1]), .G(
        dp_EBREnI2_U1_U7_clki), .Q(instr[17]) );
  LCNX1 dp_EBREnI2_U1_U0_U3 ( .CLR(n753), .D(dp_EBREnI2_m[0]), .G(
        dp_EBREnI2_U1_U7_clki), .Q(instr[16]) );
  LCNX1 dp_EBREnI3_U1_U5_U3 ( .CLR(n753), .D(dp_EBREnI3_m[5]), .G(
        dp_EBREnI3_U1_U5_clki), .Q(instr[13]) );
  LCNX1 dp_EBREnI3_U1_U4_U3 ( .CLR(n581), .D(dp_EBREnI3_m[4]), .G(
        dp_EBREnI3_U1_U5_clki), .Q(instr[12]) );
  LCNX1 dp_EBREnI3_U1_U3_U3 ( .CLR(n581), .D(dp_EBREnI3_m[3]), .G(
        dp_EBREnI3_U1_U5_clki), .Q(instr[11]) );
  LCNX1 dp_EBREnI4_U1_U7_U3 ( .CLR(n753), .D(dp_EBREnI4_m[7]), .G(
        dp_EBREnI4_U1_U7_clki), .Q(instr[7]) );
  LCNX1 dp_EBREnI4_U1_U6_U3 ( .CLR(n581), .D(dp_EBREnI4_m[6]), .G(
        dp_EBREnI4_U1_U7_clki), .Q(instr[6]) );
  LCNX1 dp_EBREnI4_U1_U5_U3 ( .CLR(n581), .D(dp_EBREnI4_m[5]), .G(
        dp_EBREnI4_U1_U7_clki), .Q(instr[5]) );
  LCNX1 dp_EBREnI4_U1_U4_U3 ( .CLR(n581), .D(dp_EBREnI4_m[4]), .G(
        dp_EBREnI4_U1_U7_clki), .Q(instr[4]) );
  LCNX1 dp_EBREnI4_U1_U3_U3 ( .CLR(n581), .D(dp_EBREnI4_m[3]), .G(
        dp_EBREnI4_U1_U7_clki), .Q(instr[3]) );
  LCNX1 dp_EBREnI4_U1_U2_U3 ( .CLR(n753), .D(dp_EBREnI4_m[2]), .G(
        dp_EBREnI4_U1_U7_clki), .Q(instr[2]) );
  LCNX1 dp_EBREnI4_U1_U1_U3 ( .CLR(n753), .D(dp_EBREnI4_m[1]), .G(
        dp_EBREnI4_U1_U7_clki), .Q(instr[1]) );
  LCX1 dp_EBL_U0_U7_U4 ( .CLR(n1), .G(dp_EBL_U0_U7_clki), .D(dp_aluresult_7_), 
        .Q(dp_EBL_m[7]) );
  LCX1 dp_EBL_U0_U6_U4 ( .CLR(n1), .G(dp_EBL_U0_U7_clki), .D(dp_aluresult_6_), 
        .Q(dp_EBL_m[6]) );
  LCX1 dp_EBL_U0_U5_U4 ( .CLR(n1), .G(dp_EBL_U0_U7_clki), .D(dp_aluresult_5_), 
        .Q(dp_EBL_m[5]) );
  LCX1 dp_EBL_U0_U4_U4 ( .CLR(n1), .G(dp_EBL_U0_U7_clki), .D(dp_aluresult_4_), 
        .Q(dp_EBL_m[4]) );
  LCX1 dp_EBL_U0_U3_U4 ( .CLR(n1), .G(dp_EBL_U0_U7_clki), .D(dp_aluresult_3_), 
        .Q(dp_EBL_m[3]) );
  LCX1 dp_EBL_U0_U2_U4 ( .CLR(n1), .G(dp_EBL_U0_U7_clki), .D(dp_aluresult_2_), 
        .Q(dp_EBL_m[2]) );
  LCX1 dp_EBL_U0_U1_U4 ( .CLR(n1), .G(dp_EBL_U0_U7_clki), .D(dp_aluresult_1_), 
        .Q(dp_EBL_m[1]) );
  LCX1 dp_EBL_U0_U0_U4 ( .CLR(n1), .G(dp_EBL_U0_U7_clki), .D(dp_aluresult_0_), 
        .Q(dp_EBL_m[0]) );
  LCX1 dp_EBB_U0_U7_U4 ( .CLR(n1), .G(dp_EBB_U0_U7_clki), .D(dp_rd2[7]), .Q(
        dp_EBB_m[7]) );
  LCX1 dp_EBB_U0_U6_U4 ( .CLR(n1), .G(dp_EBB_U0_U7_clki), .D(dp_rd2[6]), .Q(
        dp_EBB_m[6]) );
  LCX1 dp_EBB_U0_U5_U4 ( .CLR(n1), .G(dp_EBB_U0_U7_clki), .D(dp_rd2[5]), .Q(
        dp_EBB_m[5]) );
  LCX1 dp_EBB_U0_U4_U4 ( .CLR(n1), .G(dp_EBB_U0_U7_clki), .D(dp_rd2[4]), .Q(
        dp_EBB_m[4]) );
  LCX1 dp_EBB_U0_U3_U4 ( .CLR(n1), .G(dp_EBB_U0_U7_clki), .D(dp_rd2[3]), .Q(
        dp_EBB_m[3]) );
  LCX1 dp_EBB_U0_U2_U4 ( .CLR(n1), .G(dp_EBB_U0_U7_clki), .D(dp_rd2[2]), .Q(
        dp_EBB_m[2]) );
  LCX1 dp_EBB_U0_U1_U4 ( .CLR(n1), .G(dp_EBB_U0_U7_clki), .D(dp_rd2[1]), .Q(
        dp_EBB_m[1]) );
  LCX1 dp_EBB_U0_U0_U4 ( .CLR(n1), .G(dp_EBB_U0_U7_clki), .D(dp_rd2[0]), .Q(
        dp_EBB_m[0]) );
  LCX1 dp_EBA_U0_U7_U4 ( .CLR(n1), .G(dp_EBA_U0_U7_clki), .D(dp_rd1[7]), .Q(
        dp_EBA_m[7]) );
  LCX1 dp_EBA_U0_U6_U4 ( .CLR(n1), .G(dp_EBA_U0_U7_clki), .D(dp_rd1[6]), .Q(
        dp_EBA_m[6]) );
  LCX1 dp_EBA_U0_U5_U4 ( .CLR(n1), .G(dp_EBA_U0_U7_clki), .D(dp_rd1[5]), .Q(
        dp_EBA_m[5]) );
  LCX1 dp_EBA_U0_U4_U4 ( .CLR(n1), .G(dp_EBA_U0_U7_clki), .D(dp_rd1[4]), .Q(
        dp_EBA_m[4]) );
  LCX1 dp_EBA_U0_U3_U4 ( .CLR(n1), .G(dp_EBA_U0_U7_clki), .D(dp_rd1[3]), .Q(
        dp_EBA_m[3]) );
  LCX1 dp_EBA_U0_U2_U4 ( .CLR(n1), .G(dp_EBA_U0_U7_clki), .D(dp_rd1[2]), .Q(
        dp_EBA_m[2]) );
  LCX1 dp_EBA_U0_U1_U4 ( .CLR(n1), .G(dp_EBA_U0_U7_clki), .D(dp_rd1[1]), .Q(
        dp_EBA_m[1]) );
  LCX1 dp_EBA_U0_U0_U4 ( .CLR(n1), .G(dp_EBA_U0_U7_clki), .D(dp_rd1[0]), .Q(
        dp_EBA_m[0]) );
  LCX1 dp_EBM_U0_U7_U4 ( .CLR(n1), .G(dp_EBM_U0_U7_clki), .D(memdata[7]), .Q(
        dp_EBM_m[7]) );
  LCX1 dp_EBM_U0_U6_U4 ( .CLR(n1), .G(dp_EBM_U0_U7_clki), .D(memdata[6]), .Q(
        dp_EBM_m[6]) );
  LCX1 dp_EBM_U0_U5_U4 ( .CLR(n1), .G(dp_EBM_U0_U7_clki), .D(memdata[5]), .Q(
        dp_EBM_m[5]) );
  LCX1 dp_EBM_U0_U4_U4 ( .CLR(n1), .G(dp_EBM_U0_U7_clki), .D(memdata[4]), .Q(
        dp_EBM_m[4]) );
  LCX1 dp_EBM_U0_U3_U4 ( .CLR(n1), .G(dp_EBM_U0_U7_clki), .D(memdata[3]), .Q(
        dp_EBM_m[3]) );
  LCX1 dp_EBM_U0_U2_U4 ( .CLR(n1), .G(dp_EBM_U0_U7_clki), .D(memdata[2]), .Q(
        dp_EBM_m[2]) );
  LCX1 dp_EBM_U0_U1_U4 ( .CLR(n1), .G(dp_EBM_U0_U7_clki), .D(memdata[1]), .Q(
        dp_EBM_m[1]) );
  LCNX1 dp_EBL_U1_U7_U3 ( .CLR(n1), .D(dp_EBL_m[7]), .G(dp_EBL_U1_U7_clki), 
        .Q(dp_aluout_7_) );
  LCNX1 dp_EBL_U1_U6_U3 ( .CLR(n1), .D(dp_EBL_m[6]), .G(dp_EBL_U1_U7_clki), 
        .Q(dp_aluout_6_) );
  LCNX1 dp_EBL_U1_U5_U3 ( .CLR(n1), .D(dp_EBL_m[5]), .G(dp_EBL_U1_U7_clki), 
        .Q(dp_aluout_5_) );
  LCNX1 dp_EBL_U1_U4_U3 ( .CLR(n1), .D(dp_EBL_m[4]), .G(dp_EBL_U1_U7_clki), 
        .Q(dp_aluout_4_) );
  LCNX1 dp_EBL_U1_U3_U3 ( .CLR(n1), .D(dp_EBL_m[3]), .G(dp_EBL_U1_U7_clki), 
        .Q(dp_aluout_3_) );
  LCNX1 dp_EBL_U1_U2_U3 ( .CLR(n1), .D(dp_EBL_m[2]), .G(dp_EBL_U1_U7_clki), 
        .Q(dp_aluout_2_) );
  LCNX1 dp_EBL_U1_U1_U3 ( .CLR(n1), .D(dp_EBL_m[1]), .G(dp_EBL_U1_U7_clki), 
        .Q(dp_aluout_1_) );
  LCNX1 dp_EBL_U1_U0_U3 ( .CLR(n1), .D(dp_EBL_m[0]), .G(dp_EBL_U1_U7_clki), 
        .Q(dp_aluout_0_) );
  LCNX1 dp_EBB_U1_U7_U3 ( .CLR(n1), .D(dp_EBB_m[7]), .G(dp_EBB_U1_U7_clki), 
        .Q(writedata[7]) );
  LCNX1 dp_EBB_U1_U6_U3 ( .CLR(n1), .D(dp_EBB_m[6]), .G(dp_EBB_U1_U7_clki), 
        .Q(writedata[6]) );
  LCNX1 dp_EBB_U1_U5_U3 ( .CLR(n1), .D(dp_EBB_m[5]), .G(dp_EBB_U1_U7_clki), 
        .Q(writedata[5]) );
  LCNX1 dp_EBB_U1_U4_U3 ( .CLR(n1), .D(dp_EBB_m[4]), .G(dp_EBB_U1_U7_clki), 
        .Q(writedata[4]) );
  LCNX1 dp_EBB_U1_U3_U3 ( .CLR(n1), .D(dp_EBB_m[3]), .G(dp_EBB_U1_U7_clki), 
        .Q(writedata[3]) );
  LCNX1 dp_EBB_U1_U2_U3 ( .CLR(n1), .D(dp_EBB_m[2]), .G(dp_EBB_U1_U7_clki), 
        .Q(writedata[2]) );
  LCNX1 dp_EBB_U1_U1_U3 ( .CLR(n1), .D(dp_EBB_m[1]), .G(dp_EBB_U1_U7_clki), 
        .Q(writedata[1]) );
  LCNX1 dp_EBB_U1_U0_U3 ( .CLR(n1), .D(dp_EBB_m[0]), .G(dp_EBB_U1_U7_clki), 
        .Q(writedata[0]) );
  LCNX1 dp_EBA_U1_U7_U3 ( .CLR(n1), .D(dp_EBA_m[7]), .G(dp_EBA_U1_U7_clki), 
        .Q(dp_a[7]) );
  LCNX1 dp_EBA_U1_U6_U3 ( .CLR(n1), .D(dp_EBA_m[6]), .G(dp_EBA_U1_U7_clki), 
        .Q(dp_a[6]) );
  LCNX1 dp_EBA_U1_U5_U3 ( .CLR(n1), .D(dp_EBA_m[5]), .G(dp_EBA_U1_U7_clki), 
        .Q(dp_a[5]) );
  LCNX1 dp_EBA_U1_U4_U3 ( .CLR(n1), .D(dp_EBA_m[4]), .G(dp_EBA_U1_U7_clki), 
        .Q(dp_a[4]) );
  LCNX1 dp_EBA_U1_U3_U3 ( .CLR(n1), .D(dp_EBA_m[3]), .G(dp_EBA_U1_U7_clki), 
        .Q(dp_a[3]) );
  LCNX1 dp_EBA_U1_U2_U3 ( .CLR(n1), .D(dp_EBA_m[2]), .G(dp_EBA_U1_U7_clki), 
        .Q(dp_a[2]) );
  LCNX1 dp_EBA_U1_U1_U3 ( .CLR(n1), .D(dp_EBA_m[1]), .G(dp_EBA_U1_U7_clki), 
        .Q(dp_a[1]) );
  LCNX1 dp_EBA_U1_U0_U3 ( .CLR(n1), .D(dp_EBA_m[0]), .G(dp_EBA_U1_U7_clki), 
        .Q(dp_a[0]) );
  LCNX1 dp_EBM_U1_U7_U3 ( .CLR(n1), .D(dp_EBM_m[7]), .G(dp_EBM_U1_U7_clki), 
        .Q(dp_md[7]) );
  LCNX1 dp_EBM_U1_U6_U3 ( .CLR(n1), .D(dp_EBM_m[6]), .G(dp_EBM_U1_U7_clki), 
        .Q(dp_md[6]) );
  LCNX1 dp_EBM_U1_U5_U3 ( .CLR(n1), .D(dp_EBM_m[5]), .G(dp_EBM_U1_U7_clki), 
        .Q(dp_md[5]) );
  LCNX1 dp_EBM_U1_U4_U3 ( .CLR(n1), .D(dp_EBM_m[4]), .G(dp_EBM_U1_U7_clki), 
        .Q(dp_md[4]) );
  LCNX1 dp_EBM_U1_U3_U3 ( .CLR(n1), .D(dp_EBM_m[3]), .G(dp_EBM_U1_U7_clki), 
        .Q(dp_md[3]) );
  LCNX1 dp_EBM_U1_U2_U3 ( .CLR(n1), .D(dp_EBM_m[2]), .G(dp_EBM_U1_U7_clki), 
        .Q(dp_md[2]) );
  LCNX1 dp_EBM_U1_U1_U3 ( .CLR(n1), .D(dp_EBM_m[1]), .G(dp_EBM_U1_U7_clki), 
        .Q(dp_md[1]) );
  LCX1 dp_FL_EFork22_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FL_EFork22_pDFFS0_U1_di), .Q(dp_FL_EFork22_c) );
  LCX1 dp_FL_EFork22_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FL_EFork22_pDFFS1_U1_di), .Q(dp_FL_EFork22_e) );
  LCX1 dp_FL_EFork21_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FL_EFork21_pDFFS0_U1_di), .Q(dp_FL_EFork21_c) );
  LCX1 dp_FL_EFork21_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FL_EFork21_pDFFS1_U1_di), .Q(dp_FL_EFork21_e) );
  LCX1 dp_FCX_EFork21_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FCX_EFork21_pDFFS0_U1_di), .Q(dp_FCX_EFork21_c) );
  LCX1 dp_FCX_EFork21_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FCX_EFork21_pDFFS1_U1_di), .Q(dp_FCX_EFork21_e) );
  LCX1 dp_FC_EFork21_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FC_EFork21_pDFFS0_U1_di), .Q(dp_FC_EFork21_c) );
  LCX1 dp_FC_EFork21_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FC_EFork21_pDFFS1_U1_di), .Q(dp_FC_EFork21_e) );
  LCNX1 dp_FL_EFork22_pDFFS0_U0_U1 ( .CLR(n581), .D(n125), .G(clk), .Q(
        dp_FL_EFork22_pDFFS0_qi) );
  LCNX1 dp_FL_EFork22_pDFFS1_U0_U1 ( .CLR(n581), .D(dp_FL_EFork22_d), .G(clk), 
        .Q(dp_FL_EFork22_pDFFS1_qi) );
  LCNX1 dp_FL_EFork21_pDFFS0_U0_U1 ( .CLR(n753), .D(dp_FL_EFork21_b), .G(clk), 
        .Q(dp_FL_EFork21_pDFFS0_qi) );
  LCNX1 dp_FL_EFork21_pDFFS1_U0_U1 ( .CLR(n581), .D(n77), .G(clk), .Q(
        dp_FL_EFork21_pDFFS1_qi) );
  LCNX1 dp_FCX_EFork21_pDFFS0_U0_U1 ( .CLR(n581), .D(dp_FCX_EFork21_b), .G(clk), .Q(dp_FCX_EFork21_pDFFS0_qi) );
  LCNX1 dp_FCX_EFork21_pDFFS1_U0_U1 ( .CLR(n581), .D(dp_FCX_EFork21_d), .G(clk), .Q(dp_FCX_EFork21_pDFFS1_qi) );
  LCNX1 dp_FC_EFork21_pDFFS0_U0_U1 ( .CLR(n753), .D(dp_FC_EFork21_b), .G(clk), 
        .Q(dp_FC_EFork21_pDFFS0_qi) );
  LCNX1 dp_FC_EFork21_pDFFS1_U0_U1 ( .CLR(n752), .D(dp_FC_EFork21_d), .G(clk), 
        .Q(dp_FC_EFork21_pDFFS1_qi) );
  LCX1 dp_FCX_EFork31_EFork22_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FCX_EFork31_EFork22_pDFFS0_U1_di), .Q(dp_FCX_EFork31_EFork22_c) );
  LCX1 dp_FCX_EFork31_EFork22_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FCX_EFork31_EFork22_pDFFS1_U1_di), .Q(dp_FCX_EFork31_EFork22_e) );
  LCX1 dp_FCX_EFork31_EFork21_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FCX_EFork31_EFork21_pDFFS0_U1_di), .Q(dp_FCX_EFork31_EFork21_c) );
  LCX1 dp_FCX_EFork31_EFork21_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FCX_EFork31_EFork21_pDFFS1_U1_di), .Q(dp_FCX_EFork31_EFork21_e) );
  LCX1 dp_FC_EFork31_EFork22_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FC_EFork31_EFork22_pDFFS0_U1_di), .Q(dp_FC_EFork31_EFork22_c) );
  LCX1 dp_FC_EFork31_EFork22_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FC_EFork31_EFork22_pDFFS1_U1_di), .Q(dp_FC_EFork31_EFork22_e) );
  LCX1 dp_FC_EFork31_EFork21_pDFFS0_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FC_EFork31_EFork21_pDFFS0_U1_di), .Q(dp_FC_EFork31_EFork21_c) );
  LCX1 dp_FC_EFork31_EFork21_pDFFS1_U1_U3 ( .CLR(n1), .G(clk), .D(
        dp_FC_EFork31_EFork21_pDFFS1_U1_di), .Q(dp_FC_EFork31_EFork21_e) );
  LCNX1 dp_FCX_EFork31_EFork22_pDFFS0_U0_U1 ( .CLR(n753), .D(
        dp_FCX_EFork31_EFork22_b), .G(clk), .Q(
        dp_FCX_EFork31_EFork22_pDFFS0_qi) );
  LCNX1 dp_FCX_EFork31_EFork22_pDFFS1_U0_U1 ( .CLR(n581), .D(
        dp_FCX_EFork31_EFork22_d), .G(clk), .Q(
        dp_FCX_EFork31_EFork22_pDFFS1_qi) );
  LCNX1 dp_FCX_EFork31_EFork21_pDFFS0_U0_U1 ( .CLR(n581), .D(
        dp_FCX_EFork31_EFork21_b), .G(clk), .Q(
        dp_FCX_EFork31_EFork21_pDFFS0_qi) );
  LCNX1 dp_FCX_EFork31_EFork21_pDFFS1_U0_U1 ( .CLR(n753), .D(
        dp_FCX_EFork31_EFork21_d), .G(clk), .Q(
        dp_FCX_EFork31_EFork21_pDFFS1_qi) );
  LCNX1 dp_FC_EFork31_EFork22_pDFFS0_U0_U1 ( .CLR(n753), .D(
        dp_FC_EFork31_EFork22_b), .G(clk), .Q(dp_FC_EFork31_EFork22_pDFFS0_qi)
         );
  LCNX1 dp_FC_EFork31_EFork22_pDFFS1_U0_U1 ( .CLR(n581), .D(
        dp_FC_EFork31_EFork22_d), .G(clk), .Q(dp_FC_EFork31_EFork22_pDFFS1_qi)
         );
  LCNX1 dp_FC_EFork31_EFork21_pDFFS0_U0_U1 ( .CLR(n581), .D(n70), .G(clk), .Q(
        dp_FC_EFork31_EFork21_pDFFS0_qi) );
  LCNX1 dp_FC_EFork31_EFork21_pDFFS1_U0_U1 ( .CLR(n753), .D(
        dp_FC_EFork31_EFork21_d), .G(clk), .Q(dp_FC_EFork31_EFork21_pDFFS1_qi)
         );
  DCX1 dp_rfE_RAM_reg_0__0_ ( .D(n571), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_0__0_) );
  DCX1 dp_rfE_RAM_reg_0__1_ ( .D(n570), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_0__1_) );
  DCX1 dp_rfE_RAM_reg_0__2_ ( .D(n569), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_0__2_) );
  DCX1 dp_rfE_RAM_reg_0__3_ ( .D(n568), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_0__3_) );
  DCX1 dp_rfE_RAM_reg_0__4_ ( .D(n567), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_0__4_) );
  DCX1 dp_rfE_RAM_reg_0__5_ ( .D(n566), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_0__5_) );
  DCX1 dp_rfE_RAM_reg_0__6_ ( .D(n565), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_0__6_) );
  DCX1 dp_rfE_RAM_reg_0__7_ ( .D(n564), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_0__7_) );
  DCX1 dp_rfE_RAM_reg_1__0_ ( .D(n563), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_1__0_) );
  DCX1 dp_rfE_RAM_reg_1__1_ ( .D(n562), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_1__1_) );
  DCX1 dp_rfE_RAM_reg_1__2_ ( .D(n561), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_1__2_) );
  DCX1 dp_rfE_RAM_reg_1__3_ ( .D(n560), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_1__3_) );
  DCX1 dp_rfE_RAM_reg_1__4_ ( .D(n559), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_1__4_) );
  DCX1 dp_rfE_RAM_reg_1__5_ ( .D(n558), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_1__5_) );
  DCX1 dp_rfE_RAM_reg_1__6_ ( .D(n557), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_1__6_) );
  DCX1 dp_rfE_RAM_reg_1__7_ ( .D(n556), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_1__7_) );
  DCX1 dp_rfE_RAM_reg_2__0_ ( .D(n555), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_2__0_) );
  DCX1 dp_rfE_RAM_reg_2__1_ ( .D(n554), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_2__1_) );
  DCX1 dp_rfE_RAM_reg_2__2_ ( .D(n553), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_2__2_) );
  DCX1 dp_rfE_RAM_reg_2__3_ ( .D(n552), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_2__3_) );
  DCX1 dp_rfE_RAM_reg_2__4_ ( .D(n551), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_2__4_) );
  DCX1 dp_rfE_RAM_reg_2__5_ ( .D(n550), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_2__5_) );
  DCX1 dp_rfE_RAM_reg_2__6_ ( .D(n549), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_2__6_) );
  DCX1 dp_rfE_RAM_reg_2__7_ ( .D(n548), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_2__7_) );
  DCX1 dp_rfE_RAM_reg_3__0_ ( .D(n547), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_3__0_) );
  DCX1 dp_rfE_RAM_reg_3__1_ ( .D(n546), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_3__1_) );
  DCX1 dp_rfE_RAM_reg_3__2_ ( .D(n545), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_3__2_) );
  DCX1 dp_rfE_RAM_reg_3__3_ ( .D(n544), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_3__3_) );
  DCX1 dp_rfE_RAM_reg_3__4_ ( .D(n543), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_3__4_) );
  DCX1 dp_rfE_RAM_reg_3__5_ ( .D(n542), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_3__5_) );
  DCX1 dp_rfE_RAM_reg_3__6_ ( .D(n541), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_3__6_) );
  DCX1 dp_rfE_RAM_reg_3__7_ ( .D(n540), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_3__7_) );
  DCX1 dp_rfE_RAM_reg_4__0_ ( .D(n539), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_4__0_) );
  DCX1 dp_rfE_RAM_reg_4__1_ ( .D(n538), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_4__1_) );
  DCX1 dp_rfE_RAM_reg_4__2_ ( .D(n537), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_4__2_) );
  DCX1 dp_rfE_RAM_reg_4__3_ ( .D(n536), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_4__3_) );
  DCX1 dp_rfE_RAM_reg_4__4_ ( .D(n535), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_4__4_) );
  DCX1 dp_rfE_RAM_reg_4__5_ ( .D(n534), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_4__5_) );
  DCX1 dp_rfE_RAM_reg_4__6_ ( .D(n533), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_4__6_) );
  DCX1 dp_rfE_RAM_reg_4__7_ ( .D(n532), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_4__7_) );
  DCX1 dp_rfE_RAM_reg_5__0_ ( .D(n531), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_5__0_) );
  DCX1 dp_rfE_RAM_reg_5__1_ ( .D(n530), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_5__1_) );
  DCX1 dp_rfE_RAM_reg_5__2_ ( .D(n529), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_5__2_) );
  DCX1 dp_rfE_RAM_reg_5__3_ ( .D(n528), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_5__3_) );
  DCX1 dp_rfE_RAM_reg_5__4_ ( .D(n527), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_5__4_) );
  DCX1 dp_rfE_RAM_reg_5__5_ ( .D(n526), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_5__5_) );
  DCX1 dp_rfE_RAM_reg_5__6_ ( .D(n525), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_5__6_) );
  DCX1 dp_rfE_RAM_reg_5__7_ ( .D(n524), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_5__7_) );
  DCX1 dp_rfE_RAM_reg_6__0_ ( .D(n523), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_6__0_) );
  DCX1 dp_rfE_RAM_reg_6__1_ ( .D(n522), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_6__1_) );
  DCX1 dp_rfE_RAM_reg_6__2_ ( .D(n521), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_6__2_) );
  DCX1 dp_rfE_RAM_reg_6__3_ ( .D(n520), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_6__3_) );
  DCX1 dp_rfE_RAM_reg_6__4_ ( .D(n519), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_6__4_) );
  DCX1 dp_rfE_RAM_reg_6__5_ ( .D(n518), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_6__5_) );
  DCX1 dp_rfE_RAM_reg_6__6_ ( .D(n517), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_6__6_) );
  DCX1 dp_rfE_RAM_reg_6__7_ ( .D(n516), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_6__7_) );
  DCX1 dp_rfE_RAM_reg_7__0_ ( .D(n515), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_7__0_) );
  DCX1 dp_rfE_RAM_reg_7__1_ ( .D(n514), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_7__1_) );
  DCX1 dp_rfE_RAM_reg_7__2_ ( .D(n513), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_7__2_) );
  DCX1 dp_rfE_RAM_reg_7__3_ ( .D(n512), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_7__3_) );
  DCX1 dp_rfE_RAM_reg_7__4_ ( .D(n511), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_7__4_) );
  DCX1 dp_rfE_RAM_reg_7__5_ ( .D(n510), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_7__5_) );
  DCX1 dp_rfE_RAM_reg_7__6_ ( .D(n509), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_7__6_) );
  DCX1 dp_rfE_RAM_reg_7__7_ ( .D(n508), .CLK(clk), .CLR(n1), .Q(
        dp_rfE_RAM_7__7_) );
  INVX2 U123 ( .A(n378), .Y(n123) );
  OAI21X1 U192 ( .A(n589), .B(n194), .C(n195), .Y(n508) );
  NAND2X1 U193 ( .A(dp_rfE_RAM_7__7_), .B(n194), .Y(n195) );
  OAI21X1 U194 ( .A(n588), .B(n194), .C(n197), .Y(n509) );
  NAND2X1 U195 ( .A(dp_rfE_RAM_7__6_), .B(n194), .Y(n197) );
  OAI21X1 U196 ( .A(n587), .B(n194), .C(n199), .Y(n510) );
  NAND2X1 U197 ( .A(dp_rfE_RAM_7__5_), .B(n194), .Y(n199) );
  OAI21X1 U198 ( .A(n586), .B(n194), .C(n201), .Y(n511) );
  NAND2X1 U199 ( .A(dp_rfE_RAM_7__4_), .B(n194), .Y(n201) );
  OAI21X1 U200 ( .A(n585), .B(n194), .C(n203), .Y(n512) );
  NAND2X1 U201 ( .A(dp_rfE_RAM_7__3_), .B(n194), .Y(n203) );
  OAI21X1 U202 ( .A(n584), .B(n194), .C(n205), .Y(n513) );
  NAND2X1 U203 ( .A(dp_rfE_RAM_7__2_), .B(n194), .Y(n205) );
  OAI21X1 U204 ( .A(n583), .B(n194), .C(n207), .Y(n514) );
  NAND2X1 U205 ( .A(dp_rfE_RAM_7__1_), .B(n194), .Y(n207) );
  OAI21X1 U206 ( .A(n582), .B(n194), .C(n209), .Y(n515) );
  NAND2X1 U207 ( .A(dp_rfE_RAM_7__0_), .B(n194), .Y(n209) );
  OAI21X1 U209 ( .A(n589), .B(n211), .C(n212), .Y(n516) );
  NAND2X1 U210 ( .A(dp_rfE_RAM_6__7_), .B(n211), .Y(n212) );
  OAI21X1 U211 ( .A(n588), .B(n211), .C(n213), .Y(n517) );
  NAND2X1 U212 ( .A(dp_rfE_RAM_6__6_), .B(n211), .Y(n213) );
  OAI21X1 U213 ( .A(n587), .B(n211), .C(n214), .Y(n518) );
  NAND2X1 U214 ( .A(dp_rfE_RAM_6__5_), .B(n211), .Y(n214) );
  OAI21X1 U215 ( .A(n586), .B(n211), .C(n215), .Y(n519) );
  NAND2X1 U216 ( .A(dp_rfE_RAM_6__4_), .B(n211), .Y(n215) );
  OAI21X1 U217 ( .A(n585), .B(n211), .C(n216), .Y(n520) );
  NAND2X1 U218 ( .A(dp_rfE_RAM_6__3_), .B(n211), .Y(n216) );
  OAI21X1 U219 ( .A(n584), .B(n211), .C(n217), .Y(n521) );
  NAND2X1 U220 ( .A(dp_rfE_RAM_6__2_), .B(n211), .Y(n217) );
  OAI21X1 U221 ( .A(n583), .B(n211), .C(n218), .Y(n522) );
  NAND2X1 U222 ( .A(dp_rfE_RAM_6__1_), .B(n211), .Y(n218) );
  OAI21X1 U223 ( .A(n582), .B(n211), .C(n219), .Y(n523) );
  NAND2X1 U224 ( .A(dp_rfE_RAM_6__0_), .B(n211), .Y(n219) );
  NOR3X1 U226 ( .A(n96), .B(n221), .C(n222), .Y(n210) );
  OAI21X1 U227 ( .A(n589), .B(n223), .C(n224), .Y(n524) );
  NAND2X1 U228 ( .A(dp_rfE_RAM_5__7_), .B(n223), .Y(n224) );
  OAI21X1 U229 ( .A(n588), .B(n223), .C(n225), .Y(n525) );
  NAND2X1 U230 ( .A(dp_rfE_RAM_5__6_), .B(n223), .Y(n225) );
  OAI21X1 U231 ( .A(n587), .B(n223), .C(n226), .Y(n526) );
  NAND2X1 U232 ( .A(dp_rfE_RAM_5__5_), .B(n223), .Y(n226) );
  OAI21X1 U233 ( .A(n586), .B(n223), .C(n227), .Y(n527) );
  NAND2X1 U234 ( .A(dp_rfE_RAM_5__4_), .B(n223), .Y(n227) );
  OAI21X1 U235 ( .A(n585), .B(n223), .C(n228), .Y(n528) );
  NAND2X1 U236 ( .A(dp_rfE_RAM_5__3_), .B(n223), .Y(n228) );
  OAI21X1 U237 ( .A(n584), .B(n223), .C(n229), .Y(n529) );
  NAND2X1 U238 ( .A(dp_rfE_RAM_5__2_), .B(n223), .Y(n229) );
  OAI21X1 U239 ( .A(n583), .B(n223), .C(n230), .Y(n530) );
  NAND2X1 U240 ( .A(dp_rfE_RAM_5__1_), .B(n223), .Y(n230) );
  OAI21X1 U241 ( .A(n582), .B(n223), .C(n231), .Y(n531) );
  NAND2X1 U242 ( .A(dp_rfE_RAM_5__0_), .B(n223), .Y(n231) );
  OAI21X1 U244 ( .A(n589), .B(n233), .C(n234), .Y(n532) );
  NAND2X1 U245 ( .A(dp_rfE_RAM_4__7_), .B(n233), .Y(n234) );
  OAI21X1 U246 ( .A(n588), .B(n233), .C(n235), .Y(n533) );
  NAND2X1 U247 ( .A(dp_rfE_RAM_4__6_), .B(n233), .Y(n235) );
  OAI21X1 U248 ( .A(n587), .B(n233), .C(n236), .Y(n534) );
  NAND2X1 U249 ( .A(dp_rfE_RAM_4__5_), .B(n233), .Y(n236) );
  OAI21X1 U250 ( .A(n586), .B(n233), .C(n237), .Y(n535) );
  NAND2X1 U251 ( .A(dp_rfE_RAM_4__4_), .B(n233), .Y(n237) );
  OAI21X1 U252 ( .A(n585), .B(n233), .C(n238), .Y(n536) );
  NAND2X1 U253 ( .A(dp_rfE_RAM_4__3_), .B(n233), .Y(n238) );
  OAI21X1 U254 ( .A(n584), .B(n233), .C(n239), .Y(n537) );
  NAND2X1 U255 ( .A(dp_rfE_RAM_4__2_), .B(n233), .Y(n239) );
  OAI21X1 U256 ( .A(n583), .B(n233), .C(n240), .Y(n538) );
  NAND2X1 U257 ( .A(dp_rfE_RAM_4__1_), .B(n233), .Y(n240) );
  OAI21X1 U258 ( .A(n582), .B(n233), .C(n241), .Y(n539) );
  NAND2X1 U259 ( .A(dp_rfE_RAM_4__0_), .B(n233), .Y(n241) );
  NOR2X1 U261 ( .A(n222), .B(n242), .Y(n232) );
  NAND2X1 U262 ( .A(n243), .B(n221), .Y(n242) );
  OAI21X1 U263 ( .A(n589), .B(n244), .C(n245), .Y(n540) );
  NAND2X1 U264 ( .A(dp_rfE_RAM_3__7_), .B(n244), .Y(n245) );
  OAI21X1 U265 ( .A(n588), .B(n244), .C(n246), .Y(n541) );
  NAND2X1 U266 ( .A(dp_rfE_RAM_3__6_), .B(n244), .Y(n246) );
  OAI21X1 U267 ( .A(n587), .B(n244), .C(n247), .Y(n542) );
  NAND2X1 U268 ( .A(dp_rfE_RAM_3__5_), .B(n244), .Y(n247) );
  OAI21X1 U269 ( .A(n586), .B(n244), .C(n248), .Y(n543) );
  NAND2X1 U270 ( .A(dp_rfE_RAM_3__4_), .B(n244), .Y(n248) );
  OAI21X1 U271 ( .A(n585), .B(n244), .C(n249), .Y(n544) );
  NAND2X1 U272 ( .A(dp_rfE_RAM_3__3_), .B(n244), .Y(n249) );
  OAI21X1 U273 ( .A(n584), .B(n244), .C(n250), .Y(n545) );
  NAND2X1 U274 ( .A(dp_rfE_RAM_3__2_), .B(n244), .Y(n250) );
  OAI21X1 U275 ( .A(n583), .B(n244), .C(n251), .Y(n546) );
  NAND2X1 U276 ( .A(dp_rfE_RAM_3__1_), .B(n244), .Y(n251) );
  OAI21X1 U277 ( .A(n582), .B(n244), .C(n252), .Y(n547) );
  NAND2X1 U278 ( .A(dp_rfE_RAM_3__0_), .B(n244), .Y(n252) );
  OAI21X1 U280 ( .A(n589), .B(n254), .C(n255), .Y(n548) );
  NAND2X1 U281 ( .A(dp_rfE_RAM_2__7_), .B(n254), .Y(n255) );
  OAI21X1 U282 ( .A(n588), .B(n254), .C(n256), .Y(n549) );
  NAND2X1 U283 ( .A(dp_rfE_RAM_2__6_), .B(n254), .Y(n256) );
  OAI21X1 U284 ( .A(n587), .B(n254), .C(n257), .Y(n550) );
  NAND2X1 U285 ( .A(dp_rfE_RAM_2__5_), .B(n254), .Y(n257) );
  OAI21X1 U286 ( .A(n586), .B(n254), .C(n258), .Y(n551) );
  NAND2X1 U287 ( .A(dp_rfE_RAM_2__4_), .B(n254), .Y(n258) );
  OAI21X1 U288 ( .A(n585), .B(n254), .C(n259), .Y(n552) );
  NAND2X1 U289 ( .A(dp_rfE_RAM_2__3_), .B(n254), .Y(n259) );
  OAI21X1 U290 ( .A(n584), .B(n254), .C(n260), .Y(n553) );
  NAND2X1 U291 ( .A(dp_rfE_RAM_2__2_), .B(n254), .Y(n260) );
  OAI21X1 U292 ( .A(n583), .B(n254), .C(n261), .Y(n554) );
  NAND2X1 U293 ( .A(dp_rfE_RAM_2__1_), .B(n254), .Y(n261) );
  OAI21X1 U294 ( .A(n582), .B(n254), .C(n262), .Y(n555) );
  NAND2X1 U295 ( .A(dp_rfE_RAM_2__0_), .B(n254), .Y(n262) );
  NOR2X1 U297 ( .A(n221), .B(n263), .Y(n253) );
  NAND2X1 U298 ( .A(n243), .B(n222), .Y(n263) );
  OAI21X1 U299 ( .A(n589), .B(n264), .C(n265), .Y(n556) );
  NAND2X1 U300 ( .A(dp_rfE_RAM_1__7_), .B(n264), .Y(n265) );
  OAI21X1 U301 ( .A(n588), .B(n264), .C(n266), .Y(n557) );
  NAND2X1 U302 ( .A(dp_rfE_RAM_1__6_), .B(n264), .Y(n266) );
  OAI21X1 U303 ( .A(n587), .B(n264), .C(n267), .Y(n558) );
  NAND2X1 U304 ( .A(dp_rfE_RAM_1__5_), .B(n264), .Y(n267) );
  OAI21X1 U305 ( .A(n586), .B(n264), .C(n268), .Y(n559) );
  NAND2X1 U306 ( .A(dp_rfE_RAM_1__4_), .B(n264), .Y(n268) );
  OAI21X1 U307 ( .A(n585), .B(n264), .C(n269), .Y(n560) );
  NAND2X1 U308 ( .A(dp_rfE_RAM_1__3_), .B(n264), .Y(n269) );
  OAI21X1 U309 ( .A(n584), .B(n264), .C(n270), .Y(n561) );
  NAND2X1 U310 ( .A(dp_rfE_RAM_1__2_), .B(n264), .Y(n270) );
  OAI21X1 U311 ( .A(n583), .B(n264), .C(n271), .Y(n562) );
  NAND2X1 U312 ( .A(dp_rfE_RAM_1__1_), .B(n264), .Y(n271) );
  OAI21X1 U313 ( .A(n582), .B(n264), .C(n272), .Y(n563) );
  NAND2X1 U314 ( .A(dp_rfE_RAM_1__0_), .B(n264), .Y(n272) );
  OAI21X1 U316 ( .A(n589), .B(n274), .C(n275), .Y(n564) );
  NAND2X1 U317 ( .A(dp_rfE_RAM_0__7_), .B(n274), .Y(n275) );
  AOI22X1 U318 ( .A(n276), .B(dp_md[7]), .C(dp_aluout_7_), .D(n108), .Y(n193)
         );
  OAI21X1 U319 ( .A(n588), .B(n274), .C(n277), .Y(n565) );
  NAND2X1 U320 ( .A(dp_rfE_RAM_0__6_), .B(n274), .Y(n277) );
  AOI22X1 U321 ( .A(n276), .B(dp_md[6]), .C(dp_aluout_6_), .D(n108), .Y(n196)
         );
  OAI21X1 U322 ( .A(n587), .B(n274), .C(n278), .Y(n566) );
  NAND2X1 U323 ( .A(dp_rfE_RAM_0__5_), .B(n274), .Y(n278) );
  AOI22X1 U324 ( .A(n276), .B(dp_md[5]), .C(dp_aluout_5_), .D(n108), .Y(n198)
         );
  OAI21X1 U325 ( .A(n586), .B(n274), .C(n279), .Y(n567) );
  NAND2X1 U326 ( .A(dp_rfE_RAM_0__4_), .B(n274), .Y(n279) );
  AOI22X1 U327 ( .A(n276), .B(dp_md[4]), .C(dp_aluout_4_), .D(n108), .Y(n200)
         );
  OAI21X1 U328 ( .A(n585), .B(n274), .C(n280), .Y(n568) );
  NAND2X1 U329 ( .A(dp_rfE_RAM_0__3_), .B(n274), .Y(n280) );
  AOI22X1 U330 ( .A(n276), .B(dp_md[3]), .C(dp_aluout_3_), .D(n108), .Y(n202)
         );
  OAI21X1 U331 ( .A(n584), .B(n274), .C(n281), .Y(n569) );
  NAND2X1 U332 ( .A(dp_rfE_RAM_0__2_), .B(n274), .Y(n281) );
  AOI22X1 U333 ( .A(n276), .B(dp_md[2]), .C(dp_aluout_2_), .D(n108), .Y(n204)
         );
  OAI21X1 U334 ( .A(n583), .B(n274), .C(n282), .Y(n570) );
  NAND2X1 U335 ( .A(dp_rfE_RAM_0__1_), .B(n274), .Y(n282) );
  AOI22X1 U336 ( .A(n276), .B(dp_md[1]), .C(dp_aluout_1_), .D(n108), .Y(n206)
         );
  OAI21X1 U337 ( .A(n582), .B(n274), .C(n283), .Y(n571) );
  NAND2X1 U338 ( .A(dp_rfE_RAM_0__0_), .B(n274), .Y(n283) );
  NAND2X1 U341 ( .A(n222), .B(n221), .Y(n284) );
  AOI22X1 U342 ( .A(n95), .B(instr[12]), .C(instr[17]), .D(n285), .Y(n221) );
  AOI22X1 U343 ( .A(n95), .B(instr[13]), .C(instr[18]), .D(n285), .Y(n222) );
  AOI21X1 U344 ( .A(n108), .B(n285), .C(n127), .Y(n243) );
  AOI22X1 U345 ( .A(n95), .B(instr[11]), .C(instr[16]), .D(n285), .Y(n220) );
  AOI22X1 U347 ( .A(n276), .B(dp_md[0]), .C(dp_aluout_0_), .D(n108), .Y(n208)
         );
  NAND2X1 U349 ( .A(n288), .B(n289), .Y(memread) );
  NOR2X1 U350 ( .A(n290), .B(n627), .Y(dp_rd2[7]) );
  NOR2X1 U351 ( .A(n290), .B(n626), .Y(dp_rd2[6]) );
  NOR2X1 U352 ( .A(n290), .B(n625), .Y(dp_rd2[5]) );
  NOR2X1 U353 ( .A(n290), .B(n624), .Y(dp_rd2[4]) );
  NOR2X1 U354 ( .A(n290), .B(n623), .Y(dp_rd2[3]) );
  NOR2X1 U355 ( .A(n290), .B(n622), .Y(dp_rd2[2]) );
  NOR2X1 U356 ( .A(n290), .B(n621), .Y(dp_rd2[1]) );
  NOR2X1 U357 ( .A(n290), .B(n620), .Y(dp_rd2[0]) );
  NOR3X1 U358 ( .A(instr[16]), .B(instr[18]), .C(instr[17]), .Y(n290) );
  NOR2X1 U359 ( .A(n291), .B(n633), .Y(dp_rd1[7]) );
  NOR2X1 U360 ( .A(n291), .B(n632), .Y(dp_rd1[6]) );
  NOR2X1 U361 ( .A(n291), .B(n631), .Y(dp_rd1[5]) );
  NOR2X1 U362 ( .A(n291), .B(n630), .Y(dp_rd1[4]) );
  NOR2X1 U363 ( .A(n291), .B(n629), .Y(dp_rd1[3]) );
  NOR2X1 U364 ( .A(n291), .B(n628), .Y(dp_rd1[2]) );
  NOR2X1 U365 ( .A(n291), .B(n635), .Y(dp_rd1[1]) );
  NOR2X1 U366 ( .A(n291), .B(n634), .Y(dp_rd1[0]) );
  NOR3X1 U367 ( .A(instr[21]), .B(instr[23]), .C(instr[22]), .Y(n291) );
  AOI22X1 U369 ( .A(n294), .B(dp_aluout_7_), .C(n106), .D(dp_aluresult_7_), 
        .Y(n293) );
  OAI21X1 U370 ( .A(n170), .B(n292), .C(n295), .Y(dp_nextpc[6]) );
  AOI22X1 U371 ( .A(n294), .B(dp_aluout_6_), .C(n106), .D(dp_aluresult_6_), 
        .Y(n295) );
  OAI21X1 U372 ( .A(n171), .B(n292), .C(n296), .Y(dp_nextpc[5]) );
  AOI22X1 U373 ( .A(n294), .B(dp_aluout_5_), .C(n106), .D(dp_aluresult_5_), 
        .Y(n296) );
  OAI21X1 U374 ( .A(n172), .B(n292), .C(n297), .Y(dp_nextpc[4]) );
  AOI22X1 U375 ( .A(n294), .B(dp_aluout_4_), .C(n106), .D(dp_aluresult_4_), 
        .Y(n297) );
  OAI21X1 U376 ( .A(n173), .B(n292), .C(n298), .Y(dp_nextpc[3]) );
  AOI22X1 U377 ( .A(n294), .B(dp_aluout_3_), .C(n106), .D(dp_aluresult_3_), 
        .Y(n298) );
  OAI21X1 U378 ( .A(n138), .B(n292), .C(n299), .Y(dp_nextpc[2]) );
  AOI22X1 U379 ( .A(n294), .B(dp_aluout_2_), .C(n106), .D(dp_aluresult_2_), 
        .Y(n299) );
  AOI22X1 U380 ( .A(dp_aluresult_1_), .B(n106), .C(n294), .D(dp_aluout_1_), 
        .Y(n300) );
  AOI22X1 U381 ( .A(n106), .B(dp_aluresult_0_), .C(n294), .D(dp_aluout_0_), 
        .Y(n301) );
  NAND2X1 U382 ( .A(n107), .B(n292), .Y(n302) );
  MUX2NX1 U384 ( .A(DP_OP_50_64_8725_n71), .B(n105), .S(n304), .Y(
        dp_alunit_b2[6]) );
  MUX2NX1 U385 ( .A(n105), .B(DP_OP_50_64_8725_n71), .S(n305), .Y(
        dp_alunit_b2[5]) );
  MUX2NX1 U386 ( .A(DP_OP_50_64_8725_n71), .B(n105), .S(n306), .Y(
        dp_alunit_b2[4]) );
  MUX2NX1 U387 ( .A(DP_OP_50_64_8725_n71), .B(n105), .S(n307), .Y(
        dp_alunit_b2[3]) );
  MUX2NX1 U389 ( .A(DP_OP_50_64_8725_n71), .B(n105), .S(n309), .Y(
        dp_alunit_b2[1]) );
  MUX2NX1 U390 ( .A(n105), .B(DP_OP_50_64_8725_n71), .S(n310), .Y(
        dp_alunit_b2[0]) );
  NOR2X1 U391 ( .A(n161), .B(n751), .Y(dp_FX_pDFFS1_U1_di) );
  NOR2X1 U392 ( .A(n160), .B(n751), .Y(dp_FX_pDFFS0_U1_di) );
  NAND2X1 U393 ( .A(n311), .B(n312), .Y(dp_FX_d) );
  NAND2X1 U394 ( .A(n313), .B(n312), .Y(dp_FX_b) );
  OAI21X1 U395 ( .A(n67), .B(n311), .C(n313), .Y(n312) );
  NOR2X1 U396 ( .A(n155), .B(n750), .Y(dp_FP_pDFFS1_U1_di) );
  NOR2X1 U397 ( .A(n154), .B(n751), .Y(dp_FP_pDFFS0_U1_di) );
  NAND3X1 U398 ( .A(n128), .B(dp_VP), .C(n314), .Y(dp_FP_d) );
  NOR2X1 U399 ( .A(n314), .B(n128), .Y(n315) );
  NOR2X1 U400 ( .A(n175), .B(n750), .Y(dp_FL_EFork22_pDFFS1_U1_di) );
  NOR2X1 U401 ( .A(n174), .B(n751), .Y(dp_FL_EFork22_pDFFS0_U1_di) );
  NAND2X1 U402 ( .A(n126), .B(n317), .Y(dp_FL_EFork22_d) );
  NAND2X1 U403 ( .A(n318), .B(n319), .Y(n317) );
  AOI21X1 U404 ( .A(n131), .B(dp_FL_EFork22_c), .C(n320), .Y(n321) );
  NOR2X1 U405 ( .A(n177), .B(n750), .Y(dp_FL_EFork21_pDFFS1_U1_di) );
  NOR2X1 U406 ( .A(n176), .B(n750), .Y(dp_FL_EFork21_pDFFS0_U1_di) );
  NOR2X1 U407 ( .A(n320), .B(n323), .Y(n322) );
  NAND2X1 U408 ( .A(n323), .B(n320), .Y(dp_FL_EFork21_b) );
  NOR2X1 U409 ( .A(n324), .B(n325), .Y(n323) );
  NOR2X1 U410 ( .A(n185), .B(n750), .Y(dp_FCX_EFork31_EFork22_pDFFS1_U1_di) );
  NOR2X1 U411 ( .A(n184), .B(n751), .Y(dp_FCX_EFork31_EFork22_pDFFS0_U1_di) );
  NAND2X1 U412 ( .A(n326), .B(n327), .Y(dp_FCX_EFork31_EFork22_d) );
  NAND2X1 U413 ( .A(n326), .B(n328), .Y(dp_FCX_EFork31_EFork22_b) );
  NOR2X1 U414 ( .A(n146), .B(n329), .Y(n326) );
  NOR2X1 U415 ( .A(n187), .B(n750), .Y(dp_FCX_EFork31_EFork21_pDFFS1_U1_di) );
  NOR2X1 U416 ( .A(n186), .B(n750), .Y(dp_FCX_EFork31_EFork21_pDFFS0_U1_di) );
  OAI21X1 U417 ( .A(n147), .B(n183), .C(n330), .Y(dp_FCX_EFork31_EFork21_d) );
  OAI21X1 U418 ( .A(n146), .B(n182), .C(n330), .Y(dp_FCX_EFork31_EFork21_b) );
  NOR2X1 U419 ( .A(n331), .B(n74), .Y(n330) );
  NOR2X1 U420 ( .A(n179), .B(n750), .Y(dp_FCX_EFork21_pDFFS1_U1_di) );
  NOR2X1 U421 ( .A(n178), .B(n750), .Y(dp_FCX_EFork21_pDFFS0_U1_di) );
  NAND2X1 U422 ( .A(n334), .B(n335), .Y(dp_FCX_EFork21_d) );
  NAND2X1 U423 ( .A(n334), .B(n336), .Y(dp_FCX_EFork21_b) );
  NOR2X1 U424 ( .A(n147), .B(n337), .Y(n334) );
  NOR2X1 U425 ( .A(n157), .B(n750), .Y(dp_FCI2I3LM_pDFFS1_U1_di) );
  NOR2X1 U426 ( .A(n156), .B(n750), .Y(dp_FCI2I3LM_pDFFS0_U1_di) );
  NAND2X1 U427 ( .A(n339), .B(n340), .Y(dp_FCI2I3LM_d) );
  NAND2X1 U428 ( .A(dp_FCI2I3LM_e), .B(dp_SCI2I3LM2), .Y(n340) );
  NAND2X1 U429 ( .A(n339), .B(n341), .Y(dp_FCI2I3LM_b) );
  NAND2X1 U430 ( .A(dp_FCI2I3LM_c), .B(dp_SCI2I3LM1), .Y(n341) );
  NOR2X1 U431 ( .A(n342), .B(n127), .Y(n339) );
  NOR2X1 U432 ( .A(n189), .B(n749), .Y(dp_FC_EFork31_EFork22_pDFFS1_U1_di) );
  NOR2X1 U433 ( .A(n188), .B(n750), .Y(dp_FC_EFork31_EFork22_pDFFS0_U1_di) );
  NAND2X1 U434 ( .A(n343), .B(n344), .Y(dp_FC_EFork31_EFork22_d) );
  NAND2X1 U435 ( .A(n345), .B(n344), .Y(dp_FC_EFork31_EFork22_b) );
  NOR2X1 U436 ( .A(n191), .B(n749), .Y(dp_FC_EFork31_EFork21_pDFFS1_U1_di) );
  NOR2X1 U437 ( .A(n190), .B(n749), .Y(dp_FC_EFork31_EFork21_pDFFS0_U1_di) );
  NAND2X1 U438 ( .A(n71), .B(n344), .Y(dp_FC_EFork31_EFork21_d) );
  NOR2X1 U439 ( .A(n344), .B(n71), .Y(n346) );
  NOR2X1 U440 ( .A(n181), .B(n749), .Y(dp_FC_EFork21_pDFFS1_U1_di) );
  NOR2X1 U441 ( .A(n180), .B(n750), .Y(dp_FC_EFork21_pDFFS0_U1_di) );
  NAND2X1 U442 ( .A(n348), .B(n347), .Y(dp_FC_EFork21_d) );
  NAND2X1 U443 ( .A(n349), .B(n347), .Y(dp_FC_EFork21_b) );
  NOR2X1 U444 ( .A(n153), .B(n749), .Y(dp_FB_pDFFS1_U1_di) );
  NOR2X1 U445 ( .A(n152), .B(n749), .Y(dp_FB_pDFFS0_U1_di) );
  NAND2X1 U446 ( .A(n350), .B(n351), .Y(dp_FB_d) );
  NAND2X1 U447 ( .A(n352), .B(n351), .Y(dp_FB_b) );
  NOR2X1 U448 ( .A(n159), .B(n751), .Y(dp_FABCI4P_pDFFS1_U1_di) );
  NOR2X1 U449 ( .A(n158), .B(n751), .Y(dp_FABCI4P_pDFFS0_U1_di) );
  AOI21X1 U450 ( .A(dp_FABCI4P_e), .B(dp_SABCI4P2), .C(n354), .Y(n353) );
  OAI21X1 U451 ( .A(n355), .B(n143), .C(n356), .Y(dp_FABCI4P_b) );
  NOR2X1 U452 ( .A(n354), .B(n357), .Y(n356) );
  NOR2X1 U453 ( .A(n579), .B(n358), .Y(dp_EBREnP_eBCtl1_iLLS2_di) );
  AOI21X1 U454 ( .A(n314), .B(n316), .C(n145), .Y(n358) );
  NAND2X1 U455 ( .A(dp_FP_c), .B(n359), .Y(n316) );
  NAND3X1 U456 ( .A(dp_FP_e), .B(dp_VP), .C(n76), .Y(n314) );
  NOR3X1 U457 ( .A(n748), .B(dp_EBREnP_eBCtl1_b), .C(dp_EBREnP_eBCtl1_d), .Y(
        dp_EBREnP_eBCtl1_iLHS1_di) );
  NAND2X1 U458 ( .A(dp_EBREnP_eBCtl1_b), .B(dp_EBREnP_eBCtl1_d), .Y(
        dp_EBREnP_eBCtl1_f) );
  AOI21X1 U459 ( .A(n360), .B(n361), .C(dp_SABCI4LP), .Y(dp_EBREnP_eBCtl1_e)
         );
  NOR2X1 U460 ( .A(clk), .B(n362), .Y(dp_EBREnP_U0_U7_clki) );
  NAND2X1 U461 ( .A(n355), .B(pcen), .Y(n362) );
  AOI21X1 U464 ( .A(n365), .B(n366), .C(n109), .Y(n363) );
  NOR2X1 U465 ( .A(dp_aluresult_1_), .B(n738), .Y(n366) );
  OAI21X1 U467 ( .A(n739), .B(dp_src1[0]), .C(n369), .Y(n368) );
  OAI21X1 U468 ( .A(n370), .B(n371), .C(n372), .Y(n369) );
  NAND2X1 U469 ( .A(n739), .B(dp_src1[0]), .Y(n371) );
  MUX2X2 U470 ( .A(dp_pc_0_), .B(dp_a[0]), .S(n578), .Y(dp_src1[0]) );
  OAI21X1 U471 ( .A(n102), .B(n138), .C(n374), .Y(n310) );
  OAI21X1 U472 ( .A(writedata[0]), .B(n375), .C(n103), .Y(n374) );
  AOI22X1 U473 ( .A(n376), .B(dp_alunit_sum_0_), .C(n377), .D(dp_alunit_sum_7_), .Y(n367) );
  NOR2X1 U474 ( .A(n378), .B(n122), .Y(n377) );
  NAND2X1 U475 ( .A(n379), .B(n380), .Y(dp_aluresult_1_) );
  OAI21X1 U476 ( .A(n381), .B(dp_src1[1]), .C(n382), .Y(n380) );
  NOR2X1 U477 ( .A(n309), .B(n123), .Y(n382) );
  AOI22X1 U479 ( .A(n376), .B(dp_alunit_sum_1_), .C(n121), .D(dp_src1[1]), .Y(
        n379) );
  MUX2X2 U480 ( .A(dp_pc_1_), .B(dp_a[1]), .S(n618), .Y(dp_src1[1]) );
  NOR2X1 U481 ( .A(n107), .B(n385), .Y(n365) );
  NAND3X1 U482 ( .A(n386), .B(n387), .C(n388), .Y(n385) );
  NOR2X1 U483 ( .A(dp_aluresult_3_), .B(dp_aluresult_2_), .Y(n388) );
  NAND2X1 U484 ( .A(n389), .B(n390), .Y(dp_aluresult_2_) );
  OAI21X1 U485 ( .A(n381), .B(dp_src1[2]), .C(n391), .Y(n390) );
  NOR2X1 U486 ( .A(n308), .B(n123), .Y(n391) );
  OAI22X1 U488 ( .A(n393), .B(n138), .C(n102), .D(n172), .Y(n392) );
  AOI22X1 U489 ( .A(n376), .B(dp_alunit_sum_2_), .C(n121), .D(dp_src1[2]), .Y(
        n389) );
  MUX2X2 U490 ( .A(dp_pc_2_), .B(dp_a[2]), .S(n618), .Y(dp_src1[2]) );
  NAND2X1 U491 ( .A(n394), .B(n395), .Y(dp_aluresult_3_) );
  OAI21X1 U492 ( .A(n381), .B(dp_src1[3]), .C(n396), .Y(n395) );
  NOR2X1 U493 ( .A(n307), .B(n123), .Y(n396) );
  AOI21X1 U494 ( .A(n741), .B(writedata[3]), .C(n397), .Y(n307) );
  OAI22X1 U495 ( .A(n393), .B(n173), .C(n171), .D(n102), .Y(n397) );
  AOI22X1 U496 ( .A(n376), .B(dp_alunit_sum_3_), .C(n121), .D(dp_src1[3]), .Y(
        n394) );
  MUX2X2 U497 ( .A(dp_pc_3_), .B(dp_a[3]), .S(n618), .Y(dp_src1[3]) );
  NOR2X1 U498 ( .A(dp_aluresult_5_), .B(dp_aluresult_7_), .Y(n387) );
  NAND2X1 U499 ( .A(n398), .B(n399), .Y(dp_aluresult_7_) );
  OAI21X1 U500 ( .A(n381), .B(dp_src1[7]), .C(n400), .Y(n399) );
  NOR2X1 U501 ( .A(n303), .B(n123), .Y(n400) );
  AOI21X1 U502 ( .A(n741), .B(writedata[7]), .C(n401), .Y(n303) );
  OAI22X1 U503 ( .A(n393), .B(n169), .C(n102), .D(n167), .Y(n401) );
  AOI22X1 U504 ( .A(n376), .B(dp_alunit_sum_7_), .C(n121), .D(dp_src1[7]), .Y(
        n398) );
  MUX2X2 U505 ( .A(dp_pc_7_), .B(dp_a[7]), .S(n618), .Y(dp_src1[7]) );
  NAND2X1 U506 ( .A(n402), .B(n403), .Y(dp_aluresult_5_) );
  NAND2X1 U507 ( .A(n305), .B(n404), .Y(n403) );
  OAI21X1 U508 ( .A(n370), .B(n405), .C(n372), .Y(n404) );
  NAND2X1 U509 ( .A(n378), .B(n122), .Y(n370) );
  OAI21X1 U510 ( .A(n169), .B(n102), .C(n406), .Y(n305) );
  AOI22X1 U511 ( .A(n741), .B(writedata[5]), .C(n101), .D(instr[3]), .Y(n406)
         );
  AOI22X1 U512 ( .A(dp_alunit_sum_5_), .B(n376), .C(n121), .D(
        DP_OP_50_64_8725_n85), .Y(n402) );
  MUX2NX1 U513 ( .A(dp_pc_5_), .B(dp_a[5]), .S(n618), .Y(n405) );
  NOR2X1 U514 ( .A(dp_aluresult_6_), .B(dp_aluresult_4_), .Y(n386) );
  NAND2X1 U515 ( .A(n407), .B(n408), .Y(dp_aluresult_4_) );
  OAI21X1 U516 ( .A(n381), .B(dp_src1[4]), .C(n409), .Y(n408) );
  NOR2X1 U517 ( .A(n306), .B(n123), .Y(n409) );
  AOI21X1 U518 ( .A(n741), .B(writedata[4]), .C(n410), .Y(n306) );
  OAI22X1 U519 ( .A(n393), .B(n172), .C(n102), .D(n170), .Y(n410) );
  AOI22X1 U520 ( .A(n376), .B(dp_alunit_sum_4_), .C(n121), .D(dp_src1[4]), .Y(
        n407) );
  MUX2X2 U521 ( .A(dp_pc_4_), .B(dp_a[4]), .S(n618), .Y(dp_src1[4]) );
  NAND2X1 U522 ( .A(n411), .B(n412), .Y(dp_aluresult_6_) );
  OAI21X1 U523 ( .A(n381), .B(dp_src1[6]), .C(n413), .Y(n412) );
  NOR2X1 U524 ( .A(n304), .B(n123), .Y(n413) );
  AOI21X1 U525 ( .A(n741), .B(writedata[6]), .C(n414), .Y(n304) );
  OAI22X1 U526 ( .A(n393), .B(n170), .C(n102), .D(n168), .Y(n414) );
  NOR2X1 U529 ( .A(n375), .B(n415), .Y(n383) );
  OAI21X1 U532 ( .A(n418), .B(n419), .C(n744), .Y(n288) );
  AOI22X1 U533 ( .A(n376), .B(dp_alunit_sum_6_), .C(n121), .D(dp_src1[6]), .Y(
        n411) );
  MUX2X2 U534 ( .A(dp_pc_6_), .B(dp_a[6]), .S(n618), .Y(dp_src1[6]) );
  AOI21X1 U538 ( .A(n421), .B(n422), .C(n420), .Y(n378) );
  AOI21X1 U539 ( .A(instr[3]), .B(n173), .C(instr[2]), .Y(n422) );
  NOR2X1 U540 ( .A(n423), .B(instr[0]), .Y(n421) );
  AOI21X1 U541 ( .A(n424), .B(n425), .C(n420), .Y(n381) );
  AOI21X1 U542 ( .A(instr[1]), .B(instr[2]), .C(instr[0]), .Y(n425) );
  NOR2X1 U543 ( .A(dp_EBREnP_eBCtl1_b), .B(n162), .Y(dp_EBREnP_Es) );
  AOI21X1 U544 ( .A(dp_VI4), .B(n359), .C(n749), .Y(dp_EBREnI4_eBCtl1_iLLS2_di) );
  NOR3X1 U545 ( .A(n748), .B(dp_EBREnI4_eBCtl1_b), .C(dp_EBREnI4_eBCtl1_d), 
        .Y(dp_EBREnI4_eBCtl1_iLHS1_di) );
  NAND2X1 U546 ( .A(dp_EBREnI4_eBCtl1_b), .B(dp_EBREnI4_eBCtl1_d), .Y(
        dp_EBREnI4_eBCtl1_f) );
  AOI21X1 U547 ( .A(dp_FCX_EFork21_e), .B(n73), .C(dp_SCX4), .Y(
        dp_EBREnI4_eBCtl1_e) );
  NAND3X1 U548 ( .A(n426), .B(dp_EBREnI4_eBCtl1_d), .C(n427), .Y(
        dp_EBREnI4_U1_U7_clki) );
  NOR2X1 U549 ( .A(dp_EBREnI4_eBCtl1_b), .B(n65), .Y(n427) );
  NOR2X1 U550 ( .A(dp_SCX4), .B(n428), .Y(dp_EBREnI4_U0_U7_clki) );
  NAND3X1 U551 ( .A(n429), .B(n426), .C(dp_FCX_EFork21_e), .Y(n428) );
  AOI21X1 U552 ( .A(dp_VI3), .B(n319), .C(n749), .Y(dp_EBREnI3_eBCtl1_iLLS2_di) );
  NOR3X1 U553 ( .A(n748), .B(dp_EBREnI3_eBCtl1_b), .C(dp_EBREnI3_eBCtl1_d), 
        .Y(dp_EBREnI3_eBCtl1_iLHS1_di) );
  NAND2X1 U554 ( .A(dp_EBREnI3_eBCtl1_b), .B(dp_EBREnI3_eBCtl1_d), .Y(
        dp_EBREnI3_eBCtl1_f) );
  AOI21X1 U555 ( .A(dp_FCX_EFork21_c), .B(n73), .C(dp_SCX3), .Y(
        dp_EBREnI3_eBCtl1_e) );
  NAND3X1 U556 ( .A(n430), .B(dp_EBREnI3_eBCtl1_d), .C(n431), .Y(
        dp_EBREnI3_U1_U5_clki) );
  NOR2X1 U557 ( .A(dp_EBREnI3_eBCtl1_b), .B(n65), .Y(n431) );
  NOR2X1 U558 ( .A(dp_SCX3), .B(n432), .Y(dp_EBREnI3_U0_U5_clki) );
  NAND3X1 U559 ( .A(n429), .B(n430), .C(dp_FCX_EFork21_c), .Y(n432) );
  NOR2X1 U560 ( .A(clk), .B(n337), .Y(n429) );
  AOI21X1 U562 ( .A(dp_VI2), .B(n319), .C(n749), .Y(dp_EBREnI2_eBCtl1_iLLS2_di) );
  NOR3X1 U563 ( .A(n748), .B(dp_EBREnI2_eBCtl1_b), .C(dp_EBREnI2_eBCtl1_d), 
        .Y(dp_EBREnI2_eBCtl1_iLHS1_di) );
  NAND2X1 U564 ( .A(dp_EBREnI2_eBCtl1_b), .B(dp_EBREnI2_eBCtl1_d), .Y(
        dp_EBREnI2_eBCtl1_f) );
  AOI21X1 U565 ( .A(dp_FCX_EFork31_EFork22_e), .B(n72), .C(dp_SCX2), .Y(
        dp_EBREnI2_eBCtl1_e) );
  NAND3X1 U566 ( .A(n104), .B(dp_EBREnI2_eBCtl1_d), .C(n433), .Y(
        dp_EBREnI2_U1_U7_clki) );
  NOR2X1 U567 ( .A(dp_EBREnI2_eBCtl1_b), .B(n65), .Y(n433) );
  NOR2X1 U568 ( .A(dp_SCX2), .B(n434), .Y(dp_EBREnI2_U0_U7_clki) );
  NAND3X1 U569 ( .A(n435), .B(n104), .C(dp_FCX_EFork31_EFork22_e), .Y(n434) );
  NAND2X1 U570 ( .A(n419), .B(n437), .Y(n436) );
  AOI21X1 U571 ( .A(VI1), .B(n134), .C(n749), .Y(dp_EBREnI1_eBCtl1_iLLS2_di)
         );
  NOR3X1 U572 ( .A(n748), .B(dp_EBREnI1_eBCtl1_b), .C(dp_EBREnI1_eBCtl1_d), 
        .Y(dp_EBREnI1_eBCtl1_iLHS1_di) );
  NAND2X1 U573 ( .A(dp_EBREnI1_eBCtl1_b), .B(dp_EBREnI1_eBCtl1_d), .Y(
        dp_EBREnI1_eBCtl1_f) );
  AOI21X1 U574 ( .A(dp_FCX_EFork31_EFork22_c), .B(n72), .C(dp_SCX1), .Y(
        dp_EBREnI1_eBCtl1_e) );
  NAND3X1 U575 ( .A(n438), .B(dp_EBREnI1_eBCtl1_d), .C(n439), .Y(
        dp_EBREnI1_U1_U7_clki) );
  NOR2X1 U576 ( .A(dp_EBREnI1_eBCtl1_b), .B(n65), .Y(n439) );
  NOR2X1 U577 ( .A(dp_SCX1), .B(n440), .Y(dp_EBREnI1_U0_U7_clki) );
  NAND3X1 U578 ( .A(n435), .B(n438), .C(dp_FCX_EFork31_EFork22_c), .Y(n440) );
  NOR2X1 U579 ( .A(n745), .B(n441), .Y(n438) );
  NAND2X1 U580 ( .A(n418), .B(n744), .Y(n441) );
  NOR2X1 U581 ( .A(clk), .B(n329), .Y(n435) );
  NAND2X1 U582 ( .A(dp_FCX_EFork31_EFork21_c), .B(n332), .Y(n329) );
  AOI21X1 U583 ( .A(dp_VM), .B(n319), .C(n749), .Y(dp_EBM_eBCtl1_iLLS2_di) );
  NOR2X1 U584 ( .A(dp_EBM_eBCtl1_d), .B(n442), .Y(dp_EBM_eBCtl1_iLHS1_di) );
  NAND2X1 U585 ( .A(n752), .B(n151), .Y(n442) );
  NAND2X1 U586 ( .A(dp_EBM_eBCtl1_b), .B(dp_EBM_eBCtl1_d), .Y(dp_EBM_eBCtl1_f)
         );
  AOI21X1 U587 ( .A(VMemr), .B(dp_FX_e), .C(dp_SX2), .Y(dp_EBM_eBCtl1_e) );
  NAND3X1 U588 ( .A(clk), .B(dp_EBM_eBCtl1_d), .C(n151), .Y(dp_EBM_U1_U7_clki)
         );
  NOR2X1 U589 ( .A(dp_SX2), .B(n443), .Y(dp_EBM_U0_U7_clki) );
  NAND3X1 U590 ( .A(dp_FX_e), .B(VMemr), .C(n65), .Y(n443) );
  NOR2X1 U591 ( .A(n749), .B(n444), .Y(dp_EBL_eBCtl1_iLLS2_di) );
  OAI21X1 U592 ( .A(n325), .B(n324), .C(n320), .Y(n444) );
  AOI22X1 U593 ( .A(n360), .B(n131), .C(n318), .D(n319), .Y(n320) );
  NOR2X1 U594 ( .A(dp_EBL_eBCtl1_d), .B(n445), .Y(dp_EBL_eBCtl1_iLHS1_di) );
  NAND2X1 U595 ( .A(n752), .B(n148), .Y(n445) );
  NAND2X1 U596 ( .A(dp_EBL_eBCtl1_b), .B(dp_EBL_eBCtl1_d), .Y(dp_EBL_eBCtl1_f)
         );
  AOI21X1 U597 ( .A(n129), .B(dp_FABCI4P_e), .C(dp_SABCI4P2), .Y(
        dp_EBL_eBCtl1_e) );
  NAND3X1 U598 ( .A(clk), .B(dp_EBL_eBCtl1_d), .C(n148), .Y(dp_EBL_U1_U7_clki)
         );
  NOR2X1 U599 ( .A(dp_SABCI4P2), .B(n446), .Y(dp_EBL_U0_U7_clki) );
  NAND3X1 U600 ( .A(dp_FABCI4P_e), .B(n129), .C(n65), .Y(n446) );
  NOR2X1 U601 ( .A(n579), .B(n351), .Y(dp_EBB_eBCtl1_iLLS2_di) );
  AOI21X1 U602 ( .A(n352), .B(n350), .C(n144), .Y(n351) );
  NAND2X1 U603 ( .A(dp_FB_e), .B(n76), .Y(n350) );
  NAND2X1 U604 ( .A(dp_FB_c), .B(n359), .Y(n352) );
  NOR2X1 U605 ( .A(dp_EBB_eBCtl1_d), .B(n447), .Y(dp_EBB_eBCtl1_iLHS1_di) );
  NAND2X1 U606 ( .A(n752), .B(n149), .Y(n447) );
  NAND2X1 U607 ( .A(dp_EBB_eBCtl1_b), .B(dp_EBB_eBCtl1_d), .Y(dp_EBB_eBCtl1_f)
         );
  AOI21X1 U608 ( .A(n448), .B(dp_FCI2I3LM_e), .C(dp_SCI2I3LM2), .Y(
        dp_EBB_eBCtl1_e) );
  NAND3X1 U609 ( .A(clk), .B(dp_EBB_eBCtl1_d), .C(n149), .Y(dp_EBB_U1_U7_clki)
         );
  NOR2X1 U610 ( .A(dp_SCI2I3LM2), .B(n449), .Y(dp_EBB_U0_U7_clki) );
  NAND2X1 U611 ( .A(dp_FCI2I3LM_e), .B(n450), .Y(n449) );
  AOI21X1 U612 ( .A(dp_VA), .B(n359), .C(n749), .Y(dp_EBA_eBCtl1_iLLS2_di) );
  NOR2X1 U613 ( .A(dp_EBA_eBCtl1_d), .B(n451), .Y(dp_EBA_eBCtl1_iLHS1_di) );
  NAND2X1 U614 ( .A(n752), .B(n150), .Y(n451) );
  NAND2X1 U615 ( .A(dp_EBA_eBCtl1_b), .B(dp_EBA_eBCtl1_d), .Y(dp_EBA_eBCtl1_f)
         );
  AOI21X1 U616 ( .A(n448), .B(dp_FCI2I3LM_c), .C(dp_SCI2I3LM1), .Y(
        dp_EBA_eBCtl1_e) );
  NAND3X1 U617 ( .A(clk), .B(dp_EBA_eBCtl1_d), .C(n150), .Y(dp_EBA_U1_U7_clki)
         );
  NOR2X1 U618 ( .A(dp_SCI2I3LM1), .B(n452), .Y(dp_EBA_U0_U7_clki) );
  NAND2X1 U619 ( .A(dp_FCI2I3LM_c), .B(n450), .Y(n452) );
  NOR2X1 U620 ( .A(clk), .B(n127), .Y(n450) );
  NAND2X1 U621 ( .A(n453), .B(n454), .Y(cont_nextstate[3]) );
  NOR2X1 U622 ( .A(n455), .B(n456), .Y(n454) );
  AOI21X1 U623 ( .A(instr[29]), .B(n457), .C(n458), .Y(n453) );
  NAND2X1 U624 ( .A(n420), .B(n289), .Y(n458) );
  NOR2X1 U625 ( .A(n417), .B(n459), .Y(n457) );
  NAND3X1 U626 ( .A(n460), .B(n461), .C(n462), .Y(cont_nextstate[2]) );
  AOI21X1 U627 ( .A(instr[28]), .B(n456), .C(n430), .Y(n461) );
  NOR2X1 U628 ( .A(n580), .B(n463), .Y(n430) );
  NAND2X1 U629 ( .A(n619), .B(n419), .Y(n463) );
  NOR2X1 U630 ( .A(instr[27]), .B(n464), .Y(n456) );
  NAND3X1 U631 ( .A(n465), .B(n420), .C(n462), .Y(cont_nextstate[1]) );
  OAI21X1 U632 ( .A(n119), .B(n466), .C(n165), .Y(n462) );
  NOR2X1 U633 ( .A(n417), .B(instr[29]), .Y(n466) );
  AOI22X1 U634 ( .A(n467), .B(n468), .C(n437), .D(n141), .Y(n465) );
  NAND2X1 U635 ( .A(n460), .B(n469), .Y(cont_nextstate[0]) );
  AOI22X1 U636 ( .A(n165), .B(n97), .C(n419), .D(n124), .Y(n469) );
  NAND3X1 U639 ( .A(n471), .B(n467), .C(instr[31]), .Y(n459) );
  NOR2X1 U640 ( .A(instr[28]), .B(instr[27]), .Y(n467) );
  AOI21X1 U641 ( .A(instr[27]), .B(n455), .C(n426), .Y(n460) );
  NOR2X1 U642 ( .A(n580), .B(n472), .Y(n426) );
  NAND2X1 U643 ( .A(n745), .B(n418), .Y(n472) );
  NOR2X1 U644 ( .A(instr[28]), .B(n464), .Y(n455) );
  NAND2X1 U645 ( .A(n468), .B(n166), .Y(n464) );
  NOR2X1 U646 ( .A(instr[29]), .B(n473), .Y(n468) );
  NAND2X1 U647 ( .A(n119), .B(n471), .Y(n473) );
  NOR2X1 U648 ( .A(instr[26]), .B(instr[30]), .Y(n471) );
  NOR2X1 U651 ( .A(n164), .B(n751), .Y(cont_FCint_pDFFS1_U1_di) );
  NOR2X1 U652 ( .A(n163), .B(n751), .Y(cont_FCint_pDFFS0_U1_di) );
  NAND2X1 U653 ( .A(n475), .B(n476), .Y(cont_FCint_d) );
  NOR2X1 U654 ( .A(n475), .B(n476), .Y(n477) );
  NOR2X1 U655 ( .A(clk), .B(n134), .Y(cont_EBRC_lLRE1_U3_clki) );
  NAND3X1 U656 ( .A(clk), .B(cont_EBRC_eBCtl1_d), .C(n137), .Y(
        cont_EBRC_lHRE1_U3_clki) );
  NOR2X1 U657 ( .A(n476), .B(n479), .Y(cont_EBRC_eBCtl1_iLLS2_di) );
  NAND2X1 U658 ( .A(n475), .B(n581), .Y(n479) );
  NOR2X1 U659 ( .A(n344), .B(n347), .Y(n475) );
  AOI21X1 U660 ( .A(n348), .B(n349), .C(n480), .Y(n347) );
  NAND2X1 U661 ( .A(dp_FC_EFork21_c), .B(n481), .Y(n349) );
  NAND2X1 U662 ( .A(dp_FC_EFork21_e), .B(n76), .Y(n348) );
  AOI21X1 U664 ( .A(n343), .B(n345), .C(n482), .Y(n344) );
  NAND2X1 U665 ( .A(dp_FC_EFork31_EFork22_c), .B(n359), .Y(n345) );
  AOI22X1 U667 ( .A(n361), .B(n131), .C(dp_FABCI4P_e), .D(dp_SABCI4P2), .Y(
        n354) );
  AND3X1 U670 ( .A(dp_FL_EFork21_c), .B(dp_VL), .C(dp_FL_EFork22_c), .Y(n360)
         );
  NAND3X1 U672 ( .A(dp_FC_EFork31_EFork22_c), .B(dp_VB), .C(n484), .Y(n357) );
  NAND3X1 U674 ( .A(n132), .B(dp_VI4), .C(dp_FB_c), .Y(n486) );
  NAND3X1 U675 ( .A(dp_VP), .B(dp_FP_c), .C(dp_VA), .Y(n485) );
  NAND2X1 U676 ( .A(dp_FC_EFork31_EFork22_e), .B(n319), .Y(n343) );
  AOI22X1 U678 ( .A(dp_FCI2I3LM_c), .B(dp_SCI2I3LM1), .C(dp_FCI2I3LM_e), .D(
        dp_SCI2I3LM2), .Y(n342) );
  NAND3X1 U681 ( .A(cont_FCint_e), .B(cont_VCint), .C(dp_FC_EFork31_EFork21_c), 
        .Y(n482) );
  AND3X1 U683 ( .A(dp_FL_EFork21_c), .B(dp_FL_EFork22_e), .C(dp_VL), .Y(n318)
         );
  NOR2X1 U684 ( .A(n478), .B(n489), .Y(n476) );
  NAND2X1 U685 ( .A(cont_VCint), .B(cont_FCint_c), .Y(n489) );
  NOR2X1 U686 ( .A(cont_SCI1), .B(n490), .Y(n478) );
  NOR3X1 U687 ( .A(n748), .B(cont_EBRC_eBCtl1_b), .C(cont_EBRC_eBCtl1_d), .Y(
        cont_EBRC_eBCtl1_iLHS1_di) );
  NAND2X1 U689 ( .A(cont_EBRC_eBCtl1_b), .B(cont_EBRC_eBCtl1_d), .Y(
        cont_EBRC_eBCtl1_f) );
  NOR2X1 U690 ( .A(cont_SCI1), .B(n133), .Y(cont_EBRC_eBCtl1_e) );
  NAND3X1 U691 ( .A(cont_VCint), .B(cont_FCint_c), .C(VI1), .Y(n490) );
  OAI21X1 U692 ( .A(n491), .B(n420), .C(n107), .Y(alucont_2_) );
  AOI21X1 U699 ( .A(instr[0]), .B(n172), .C(n492), .Y(n491) );
  NAND2X1 U700 ( .A(n173), .B(n424), .Y(n492) );
  NOR2X1 U701 ( .A(instr[3]), .B(n423), .Y(n424) );
  NAND2X1 U702 ( .A(instr[5]), .B(n170), .Y(n423) );
  OAI22X1 U703 ( .A(n118), .B(dp_pc_7_), .C(dp_aluout_7_), .D(n494), .Y(n493)
         );
  OAI22X1 U704 ( .A(n118), .B(dp_pc_6_), .C(dp_aluout_6_), .D(n494), .Y(n495)
         );
  OAI22X1 U705 ( .A(n118), .B(dp_pc_5_), .C(dp_aluout_5_), .D(n494), .Y(n496)
         );
  OAI22X1 U706 ( .A(n118), .B(dp_pc_4_), .C(dp_aluout_4_), .D(n494), .Y(n497)
         );
  OAI22X1 U707 ( .A(n118), .B(dp_pc_3_), .C(dp_aluout_3_), .D(n494), .Y(n498)
         );
  OAI22X1 U708 ( .A(n118), .B(dp_pc_2_), .C(dp_aluout_2_), .D(n494), .Y(n499)
         );
  OAI22X1 U709 ( .A(n118), .B(dp_pc_1_), .C(dp_aluout_1_), .D(n494), .Y(n500)
         );
  OAI22X1 U710 ( .A(n118), .B(dp_pc_0_), .C(dp_aluout_0_), .D(n494), .Y(n501)
         );
  NOR3X1 U712 ( .A(n744), .B(n745), .C(n474), .Y(memwrite) );
  NAND2X1 U714 ( .A(n502), .B(n470), .Y(n289) );
  NOR2X1 U716 ( .A(n580), .B(n124), .Y(n502) );
  NAND3X1 U718 ( .A(dp_VB), .B(n136), .C(dp_FP_e), .Y(n504) );
  NAND3X1 U719 ( .A(dp_FB_e), .B(dp_FC_EFork21_e), .C(n505), .Y(n503) );
  NOR2X1 U720 ( .A(n325), .B(n145), .Y(n505) );
  NAND2X1 U721 ( .A(dp_VL), .B(dp_FL_EFork21_e), .Y(n325) );
  NAND2X1 U722 ( .A(n313), .B(n311), .Y(SMemr) );
  NAND2X1 U724 ( .A(n68), .B(n481), .Y(n313) );
  NAND2X1 U725 ( .A(n331), .B(n332), .Y(n481) );
  NAND2X1 U727 ( .A(n136), .B(dp_FC_EFork21_c), .Y(n507) );
  NAND3X1 U728 ( .A(cont_FCint_e), .B(cont_VCint), .C(dp_FC_EFork31_EFork21_e), 
        .Y(n480) );
  AOI22X1 U729 ( .A(dp_FCX_EFork31_EFork21_c), .B(n333), .C(
        dp_FCX_EFork31_EFork21_e), .D(n338), .Y(n331) );
  NAND2X1 U730 ( .A(n336), .B(n335), .Y(n338) );
  NAND2X1 U731 ( .A(dp_FCX_EFork21_e), .B(dp_SCX4), .Y(n335) );
  NAND2X1 U732 ( .A(dp_FCX_EFork21_c), .B(dp_SCX3), .Y(n336) );
  NAND2X1 U733 ( .A(n328), .B(n327), .Y(n333) );
  NAND2X1 U734 ( .A(dp_FCX_EFork31_EFork22_e), .B(dp_SCX2), .Y(n327) );
  NAND2X1 U735 ( .A(dp_FCX_EFork31_EFork22_c), .B(dp_SCX1), .Y(n328) );
  INVX1 U122 ( .A(n381), .Y(n122) );
  NOR2X2 U668 ( .A(dp_SABCI4LP), .B(n483), .Y(n355) );
  INVX1 U145 ( .A(dp_VP), .Y(n145) );
  NOR2X2 U663 ( .A(n135), .B(SMeml), .Y(n324) );
  INVX1 U126 ( .A(n320), .Y(n126) );
  INVX1 U71 ( .A(n347), .Y(n71) );
  INVX1 U100 ( .A(n300), .Y(n100) );
  INVX1 U182 ( .A(dp_FCX_EFork31_EFork21_c), .Y(n182) );
  INVX1 U74 ( .A(n332), .Y(n74) );
  INVX1 U183 ( .A(dp_FCX_EFork31_EFork21_e), .Y(n183) );
  INVX1 U166 ( .A(instr[31]), .Y(n166) );
  INVX1 U109 ( .A(n288), .Y(n109) );
  INVX1 U162 ( .A(dp_EBREnP_eBCtl1_d), .Y(n162) );
  NAND2X1 U561 ( .A(dp_FCX_EFork31_EFork21_e), .B(n332), .Y(n337) );
  INVX2 U142 ( .A(cont_state_1_), .Y(n142) );
  NAND2X1 U713 ( .A(n142), .B(n619), .Y(n474) );
  INVX2 U106 ( .A(n302), .Y(n106) );
  INVX1 U171 ( .A(instr[3]), .Y(n171) );
  INVX2 U99 ( .A(n405), .Y(DP_OP_50_64_8725_n85) );
  NAND2X1 U536 ( .A(n381), .B(n378), .Y(n372) );
  INVX2 U121 ( .A(n372), .Y(n121) );
  INVX2 U132 ( .A(n482), .Y(n132) );
  INVX2 U131 ( .A(n355), .Y(n131) );
  NAND2X2 U666 ( .A(n129), .B(n354), .Y(n359) );
  INVX2 U128 ( .A(n316), .Y(n128) );
  NOR2X2 U717 ( .A(n503), .B(n504), .Y(VMeml) );
  INVX2 U135 ( .A(VMeml), .Y(n135) );
  INVX2 U76 ( .A(n324), .Y(n76) );
  INVX1 U144 ( .A(dp_VB), .Y(n144) );
  INVX1 U148 ( .A(dp_EBL_eBCtl1_b), .Y(n148) );
  INVX1 U149 ( .A(dp_EBB_eBCtl1_b), .Y(n149) );
  INVX1 U150 ( .A(dp_EBA_eBCtl1_b), .Y(n150) );
  INVX1 U151 ( .A(dp_EBM_eBCtl1_b), .Y(n151) );
  INVX2 U127 ( .A(n448), .Y(n127) );
  NAND2X1 U723 ( .A(dp_FX_e), .B(dp_SX2), .Y(n311) );
  INVX2 U146 ( .A(n333), .Y(n146) );
  INVX2 U147 ( .A(n338), .Y(n147) );
  INVX2 U72 ( .A(n329), .Y(n72) );
  INVX2 U73 ( .A(n337), .Y(n73) );
  INVX2 U165 ( .A(n459), .Y(n165) );
  INVX2 U96 ( .A(n243), .Y(n96) );
  INVX2 U112 ( .A(n499), .Y(adr[2]) );
  INVX2 U110 ( .A(n501), .Y(adr[0]) );
  INVX2 U111 ( .A(n500), .Y(adr[1]) );
  INVX2 U117 ( .A(n493), .Y(adr[7]) );
  INVX2 U116 ( .A(n495), .Y(adr[6]) );
  INVX2 U114 ( .A(n497), .Y(adr[4]) );
  INVX2 U115 ( .A(n496), .Y(adr[5]) );
  INVX2 U113 ( .A(n498), .Y(adr[3]) );
  INVX2 U104 ( .A(n436), .Y(n104) );
  INVX1 U137 ( .A(cont_EBRC_eBCtl1_b), .Y(n137) );
  NOR2X2 U671 ( .A(n357), .B(n143), .Y(n361) );
  INVX1 U67 ( .A(VMemr), .Y(n67) );
  INVX2 U118 ( .A(n494), .Y(n118) );
  INVX2 U65 ( .A(clk), .Y(n65) );
  INVX1 U101 ( .A(n393), .Y(n101) );
  NAND2X1 U736 ( .A(VMemr), .B(dp_FX_c), .Y(n506) );
  NAND2X1 U463 ( .A(n580), .B(n364), .Y(n292) );
  NOR2X1 U537 ( .A(n381), .B(n378), .Y(n376) );
  INVX1 U129 ( .A(n357), .Y(n129) );
  NAND2X1 U346 ( .A(n619), .B(n286), .Y(n285) );
  INVX2 U103 ( .A(n415), .Y(n103) );
  NAND2X2 U669 ( .A(n360), .B(n361), .Y(n483) );
  INVX2 U108 ( .A(n276), .Y(n108) );
  NOR2X1 U340 ( .A(n96), .B(n284), .Y(n273) );
  INVX1 U119 ( .A(n416), .Y(n119) );
  NAND2X1 U315 ( .A(n273), .B(n94), .Y(n264) );
  NAND2X1 U279 ( .A(n253), .B(n94), .Y(n244) );
  NAND2X1 U243 ( .A(n232), .B(n94), .Y(n223) );
  NAND2X1 U208 ( .A(n210), .B(n94), .Y(n194) );
  INVX1 U181 ( .A(dp_FC_EFork21_pDFFS1_qi), .Y(n181) );
  INVX1 U153 ( .A(dp_FB_pDFFS1_qi), .Y(n153) );
  INVX1 U152 ( .A(dp_FB_pDFFS0_qi), .Y(n152) );
  INVX1 U159 ( .A(dp_FABCI4P_pDFFS1_qi), .Y(n159) );
  INVX1 U191 ( .A(dp_FC_EFork31_EFork21_pDFFS1_qi), .Y(n191) );
  INVX1 U157 ( .A(dp_FCI2I3LM_pDFFS1_qi), .Y(n157) );
  INVX1 U188 ( .A(dp_FC_EFork31_EFork22_pDFFS0_qi), .Y(n188) );
  INVX1 U185 ( .A(dp_FCX_EFork31_EFork22_pDFFS1_qi), .Y(n185) );
  INVX2 U143 ( .A(dp_FABCI4P_c), .Y(n143) );
  INVX1 U179 ( .A(dp_FCX_EFork21_pDFFS1_qi), .Y(n179) );
  INVX1 U189 ( .A(dp_FC_EFork31_EFork22_pDFFS1_qi), .Y(n189) );
  INVX1 U190 ( .A(dp_FC_EFork31_EFork21_pDFFS0_qi), .Y(n190) );
  INVX1 U177 ( .A(dp_FL_EFork21_pDFFS1_qi), .Y(n177) );
  INVX1 U184 ( .A(dp_FCX_EFork31_EFork22_pDFFS0_qi), .Y(n184) );
  INVX1 U158 ( .A(dp_FABCI4P_pDFFS0_qi), .Y(n158) );
  INVX1 U154 ( .A(dp_FP_pDFFS0_qi), .Y(n154) );
  INVX1 U161 ( .A(dp_FX_pDFFS1_qi), .Y(n161) );
  INVX1 U175 ( .A(dp_FL_EFork22_pDFFS1_qi), .Y(n175) );
  INVX1 U155 ( .A(dp_FP_pDFFS1_qi), .Y(n155) );
  INVX1 U164 ( .A(cont_FCint_pDFFS1_qi), .Y(n164) );
  INVX1 U174 ( .A(dp_FL_EFork22_pDFFS0_qi), .Y(n174) );
  INVX1 U178 ( .A(dp_FCX_EFork21_pDFFS0_qi), .Y(n178) );
  INVX1 U176 ( .A(dp_FL_EFork21_pDFFS0_qi), .Y(n176) );
  INVX1 U163 ( .A(cont_FCint_pDFFS0_qi), .Y(n163) );
  INVX1 U180 ( .A(dp_FC_EFork21_pDFFS0_qi), .Y(n180) );
  INVX1 U187 ( .A(dp_FCX_EFork31_EFork21_pDFFS1_qi), .Y(n187) );
  INVX1 U160 ( .A(dp_FX_pDFFS0_qi), .Y(n160) );
  INVX1 U186 ( .A(dp_FCX_EFork31_EFork21_pDFFS0_qi), .Y(n186) );
  INVX1 U156 ( .A(dp_FCI2I3LM_pDFFS0_qi), .Y(n156) );
  INVX1 U68 ( .A(n506), .Y(n68) );
  INVX1 U136 ( .A(n480), .Y(n136) );
  INVX1 U133 ( .A(n490), .Y(n133) );
  INVX1 U134 ( .A(n478), .Y(n134) );
  NOR2X1 U673 ( .A(n485), .B(n486), .Y(n484) );
  NOR2X1 U726 ( .A(n506), .B(n507), .Y(n332) );
  NOR2X1 U650 ( .A(n141), .B(n474), .Y(n364) );
  INVX1 U120 ( .A(n289), .Y(n120) );
  INVX1 U95 ( .A(n285), .Y(n95) );
  INVX1 U167 ( .A(instr[7]), .Y(n167) );
  INVX1 U168 ( .A(instr[6]), .Y(n168) );
  INVX2 U172 ( .A(instr[2]), .Y(n172) );
  INVX2 U138 ( .A(instr[0]), .Y(n138) );
  INVX2 U170 ( .A(instr[4]), .Y(n170) );
  INVX2 U173 ( .A(instr[1]), .Y(n173) );
  INVX1 U77 ( .A(n322), .Y(n77) );
  INVX1 U125 ( .A(n321), .Y(n125) );
  INVX1 U130 ( .A(n353), .Y(n130) );
  INVX1 U94 ( .A(n220), .Y(n94) );
  INVX1 U70 ( .A(n346), .Y(n70) );
  INVX1 U75 ( .A(n315), .Y(n75) );
  INVX1 U69 ( .A(n477), .Y(n69) );
  NAND2X1 U737 ( .A(n375), .B(n415), .Y(n393) );
  INVX2 U738 ( .A(n740), .Y(n741) );
  NAND2X1 U739 ( .A(n448), .B(n342), .Y(n319) );
  INVX2 U740 ( .A(cont_state_3_), .Y(n744) );
  NOR2X1 U741 ( .A(n744), .B(n140), .Y(n286) );
  NOR2X1 U742 ( .A(cont_state_1_), .B(n619), .Y(n418) );
  NOR2X1 U743 ( .A(n141), .B(n142), .Y(n470) );
  INVX1 U744 ( .A(n102), .Y(n573) );
  AOI22X1 U745 ( .A(n741), .B(writedata[1]), .C(instr[1]), .D(n573), .Y(n309)
         );
  MUX2NX1 U746 ( .A(DP_OP_50_64_8725_n71), .B(n105), .S(n303), .Y(n574) );
  XOR2X1 U747 ( .A(n574), .B(dp_src1[7]), .Y(n575) );
  XNOR2X1 U748 ( .A(n609), .B(n575), .Y(dp_alunit_sum_7_) );
  NAND3X1 U749 ( .A(n132), .B(dp_VM), .C(dp_VI2), .Y(n576) );
  NAND3X1 U750 ( .A(dp_FC_EFork31_EFork22_e), .B(n318), .C(dp_VI3), .Y(n577)
         );
  NOR2X1 U751 ( .A(n576), .B(n577), .Y(n448) );
  NAND3X1 U752 ( .A(n417), .B(n107), .C(n420), .Y(n578) );
  INVX2 U753 ( .A(n294), .Y(n107) );
  NOR2X2 U754 ( .A(n141), .B(n287), .Y(n294) );
  BUFX4 U755 ( .A(reset), .Y(n579) );
  BUFX4 U756 ( .A(alucont_2_), .Y(DP_OP_50_64_8725_n71) );
  BUFX2 U757 ( .A(n196), .Y(n588) );
  BUFX2 U758 ( .A(n208), .Y(n582) );
  BUFX2 U759 ( .A(n206), .Y(n583) );
  BUFX2 U760 ( .A(n204), .Y(n584) );
  BUFX2 U761 ( .A(n202), .Y(n585) );
  BUFX2 U762 ( .A(n200), .Y(n586) );
  BUFX2 U763 ( .A(n198), .Y(n587) );
  INVX1 U764 ( .A(n292), .Y(n746) );
  INVX4 U765 ( .A(n744), .Y(n580) );
  BUFX4 U766 ( .A(cont_state_2_), .Y(n745) );
  INVX1 U767 ( .A(writedata[2]), .Y(n742) );
  BUFX2 U768 ( .A(cont_state_0_), .Y(n619) );
  INVX4 U769 ( .A(n579), .Y(n581) );
  BUFX2 U770 ( .A(n193), .Y(n589) );
  XOR2X1 U771 ( .A(dp_src1[0]), .B(dp_alunit_b2[0]), .Y(n590) );
  XOR2X1 U772 ( .A(n613), .B(DP_OP_50_64_8725_n71), .Y(dp_alunit_sum_0_) );
  AOI22X1 U773 ( .A(dp_alunit_b2[0]), .B(dp_src1[0]), .C(DP_OP_50_64_8725_n71), 
        .D(n590), .Y(n594) );
  XOR2X1 U774 ( .A(dp_alunit_b2[1]), .B(dp_src1[1]), .Y(n591) );
  XNOR2X1 U775 ( .A(n611), .B(n591), .Y(dp_alunit_sum_1_) );
  XOR2X1 U776 ( .A(dp_alunit_b2[2]), .B(dp_src1[2]), .Y(n596) );
  NOR2X1 U777 ( .A(dp_src1[1]), .B(dp_alunit_b2[1]), .Y(n593) );
  NAND2X1 U778 ( .A(dp_src1[1]), .B(dp_alunit_b2[1]), .Y(n592) );
  OAI21X1 U779 ( .A(n594), .B(n593), .C(n592), .Y(n595) );
  XOR2X1 U780 ( .A(n616), .B(n615), .Y(dp_alunit_sum_2_) );
  AOI22X1 U781 ( .A(dp_alunit_b2[2]), .B(dp_src1[2]), .C(n596), .D(n595), .Y(
        n600) );
  XOR2X1 U782 ( .A(dp_alunit_b2[3]), .B(dp_src1[3]), .Y(n597) );
  XNOR2X1 U783 ( .A(n610), .B(n597), .Y(dp_alunit_sum_3_) );
  XOR2X1 U784 ( .A(dp_alunit_b2[4]), .B(dp_src1[4]), .Y(n602) );
  NOR2X1 U785 ( .A(dp_src1[3]), .B(dp_alunit_b2[3]), .Y(n599) );
  NAND2X1 U786 ( .A(dp_src1[3]), .B(dp_alunit_b2[3]), .Y(n598) );
  OAI21X1 U787 ( .A(n600), .B(n599), .C(n598), .Y(n601) );
  XOR2X1 U788 ( .A(n602), .B(n614), .Y(dp_alunit_sum_4_) );
  AOI22X1 U789 ( .A(dp_alunit_b2[4]), .B(dp_src1[4]), .C(n602), .D(n601), .Y(
        n606) );
  XOR2X1 U790 ( .A(dp_alunit_b2[5]), .B(DP_OP_50_64_8725_n85), .Y(n603) );
  XNOR2X1 U791 ( .A(n612), .B(n603), .Y(dp_alunit_sum_5_) );
  XOR2X1 U792 ( .A(dp_alunit_b2[6]), .B(dp_src1[6]), .Y(n608) );
  NOR2X1 U793 ( .A(DP_OP_50_64_8725_n85), .B(dp_alunit_b2[5]), .Y(n605) );
  NAND2X1 U794 ( .A(DP_OP_50_64_8725_n85), .B(dp_alunit_b2[5]), .Y(n604) );
  OAI21X1 U795 ( .A(n606), .B(n605), .C(n604), .Y(n607) );
  XOR2X1 U796 ( .A(n608), .B(n617), .Y(dp_alunit_sum_6_) );
  AOI22X1 U797 ( .A(dp_alunit_b2[6]), .B(dp_src1[6]), .C(n608), .D(n607), .Y(
        n609) );
  AOI22X1 U798 ( .A(dp_alunit_b2[2]), .B(dp_src1[2]), .C(n616), .D(n615), .Y(
        n610) );
  BUFX2 U799 ( .A(n594), .Y(n611) );
  AOI22X1 U800 ( .A(dp_alunit_b2[4]), .B(dp_src1[4]), .C(n602), .D(n614), .Y(
        n612) );
  BUFX2 U801 ( .A(n590), .Y(n613) );
  BUFX2 U802 ( .A(n601), .Y(n614) );
  BUFX2 U803 ( .A(n595), .Y(n615) );
  BUFX2 U804 ( .A(n596), .Y(n616) );
  BUFX2 U805 ( .A(n607), .Y(n617) );
  BUFX2 U806 ( .A(n578), .Y(n618) );
  NOR2X1 U807 ( .A(n580), .B(n619), .Y(n437) );
  NAND2X2 U808 ( .A(n580), .B(n418), .Y(n287) );
  NAND2X1 U809 ( .A(n220), .B(n210), .Y(n211) );
  BUFX2 U810 ( .A(instr[21]), .Y(n736) );
  BUFX2 U811 ( .A(instr[21]), .Y(n735) );
  BUFX2 U812 ( .A(instr[16]), .Y(n685) );
  BUFX2 U813 ( .A(instr[16]), .Y(n684) );
  INVX2 U814 ( .A(n579), .Y(n752) );
  NAND2X1 U815 ( .A(n220), .B(n273), .Y(n274) );
  NAND2X1 U816 ( .A(n220), .B(n232), .Y(n233) );
  NAND2X1 U817 ( .A(n220), .B(n253), .Y(n254) );
  NOR2X1 U818 ( .A(n745), .B(n287), .Y(n276) );
  BUFX2 U819 ( .A(instr[17]), .Y(n686) );
  NAND2X2 U820 ( .A(n416), .B(n417), .Y(n415) );
  NOR2X1 U821 ( .A(n120), .B(memwrite), .Y(n494) );
  BUFX2 U822 ( .A(instr[22]), .Y(n737) );
  BUFX2 U823 ( .A(reset), .Y(n749) );
  NOR2X2 U824 ( .A(n375), .B(n103), .Y(n384) );
  INVX4 U825 ( .A(n384), .Y(n102) );
  NAND2X2 U826 ( .A(n416), .B(n288), .Y(n375) );
  NAND2X2 U827 ( .A(n744), .B(n364), .Y(n416) );
  INVX4 U828 ( .A(DP_OP_50_64_8725_n71), .Y(n105) );
  INVX2 U829 ( .A(n579), .Y(n753) );
  NAND2X1 U830 ( .A(n363), .B(n292), .Y(pcen) );
  BUFX4 U831 ( .A(reset), .Y(n750) );
  NAND2X2 U832 ( .A(n437), .B(n470), .Y(n417) );
  BUFX4 U833 ( .A(reset), .Y(n751) );
  BUFX4 U834 ( .A(reset), .Y(n748) );
  INVX2 U835 ( .A(n383), .Y(n740) );
  INVX1 U836 ( .A(n619), .Y(n124) );
  INVX2 U837 ( .A(n419), .Y(n140) );
  MUX2NX1 U838 ( .A(n640), .B(n641), .S(instr[18]), .Y(n620) );
  MUX2NX1 U839 ( .A(n646), .B(n647), .S(instr[18]), .Y(n621) );
  MUX2NX1 U840 ( .A(n652), .B(n653), .S(instr[18]), .Y(n622) );
  MUX2NX1 U841 ( .A(n658), .B(n659), .S(instr[18]), .Y(n623) );
  MUX2NX1 U842 ( .A(n664), .B(n665), .S(instr[18]), .Y(n624) );
  MUX2NX1 U843 ( .A(n670), .B(n671), .S(instr[18]), .Y(n625) );
  MUX2NX1 U844 ( .A(n676), .B(n677), .S(instr[18]), .Y(n626) );
  MUX2NX1 U845 ( .A(n682), .B(n683), .S(instr[18]), .Y(n627) );
  MUX2NX1 U846 ( .A(n703), .B(n704), .S(instr[23]), .Y(n628) );
  MUX2NX1 U847 ( .A(n709), .B(n710), .S(instr[23]), .Y(n629) );
  MUX2NX1 U848 ( .A(n715), .B(n716), .S(instr[23]), .Y(n630) );
  MUX2NX1 U849 ( .A(n721), .B(n722), .S(instr[23]), .Y(n631) );
  MUX2NX1 U850 ( .A(n727), .B(n728), .S(instr[23]), .Y(n632) );
  MUX2NX1 U851 ( .A(n733), .B(n734), .S(instr[23]), .Y(n633) );
  MUX2NX1 U852 ( .A(n691), .B(n692), .S(instr[23]), .Y(n634) );
  MUX2NX1 U853 ( .A(n697), .B(n698), .S(instr[23]), .Y(n635) );
  TIEHI U854 ( .Y(n1) );
  MUX2NX1 U855 ( .A(dp_rfE_RAM_0__0_), .B(dp_rfE_RAM_1__0_), .S(n685), .Y(n636) );
  MUX2NX1 U856 ( .A(dp_rfE_RAM_2__0_), .B(dp_rfE_RAM_3__0_), .S(n685), .Y(n637) );
  MUX2NX1 U857 ( .A(dp_rfE_RAM_4__0_), .B(dp_rfE_RAM_5__0_), .S(n685), .Y(n638) );
  MUX2NX1 U858 ( .A(dp_rfE_RAM_6__0_), .B(dp_rfE_RAM_7__0_), .S(n685), .Y(n639) );
  MUX2NX1 U859 ( .A(n636), .B(n637), .S(n686), .Y(n640) );
  MUX2NX1 U860 ( .A(n638), .B(n639), .S(n686), .Y(n641) );
  MUX2NX1 U861 ( .A(dp_rfE_RAM_0__1_), .B(dp_rfE_RAM_1__1_), .S(n684), .Y(n642) );
  MUX2NX1 U862 ( .A(dp_rfE_RAM_2__1_), .B(dp_rfE_RAM_3__1_), .S(n684), .Y(n643) );
  MUX2NX1 U863 ( .A(dp_rfE_RAM_4__1_), .B(dp_rfE_RAM_5__1_), .S(n684), .Y(n644) );
  MUX2NX1 U864 ( .A(dp_rfE_RAM_6__1_), .B(dp_rfE_RAM_7__1_), .S(n684), .Y(n645) );
  MUX2NX1 U865 ( .A(n642), .B(n643), .S(n686), .Y(n646) );
  MUX2NX1 U866 ( .A(n644), .B(n645), .S(n686), .Y(n647) );
  MUX2NX1 U867 ( .A(dp_rfE_RAM_0__2_), .B(dp_rfE_RAM_1__2_), .S(n684), .Y(n648) );
  MUX2NX1 U868 ( .A(dp_rfE_RAM_2__2_), .B(dp_rfE_RAM_3__2_), .S(n684), .Y(n649) );
  MUX2NX1 U869 ( .A(dp_rfE_RAM_4__2_), .B(dp_rfE_RAM_5__2_), .S(n684), .Y(n650) );
  MUX2NX1 U870 ( .A(dp_rfE_RAM_6__2_), .B(dp_rfE_RAM_7__2_), .S(n684), .Y(n651) );
  MUX2NX1 U871 ( .A(n648), .B(n649), .S(n686), .Y(n652) );
  MUX2NX1 U872 ( .A(n650), .B(n651), .S(n686), .Y(n653) );
  MUX2NX1 U873 ( .A(dp_rfE_RAM_0__3_), .B(dp_rfE_RAM_1__3_), .S(n684), .Y(n654) );
  MUX2NX1 U874 ( .A(dp_rfE_RAM_2__3_), .B(dp_rfE_RAM_3__3_), .S(n684), .Y(n655) );
  MUX2NX1 U875 ( .A(dp_rfE_RAM_4__3_), .B(dp_rfE_RAM_5__3_), .S(n684), .Y(n656) );
  MUX2NX1 U876 ( .A(dp_rfE_RAM_6__3_), .B(dp_rfE_RAM_7__3_), .S(n684), .Y(n657) );
  MUX2NX1 U877 ( .A(n654), .B(n655), .S(n686), .Y(n658) );
  MUX2NX1 U878 ( .A(n656), .B(n657), .S(n686), .Y(n659) );
  MUX2NX1 U879 ( .A(dp_rfE_RAM_0__4_), .B(dp_rfE_RAM_1__4_), .S(n684), .Y(n660) );
  MUX2NX1 U880 ( .A(dp_rfE_RAM_2__4_), .B(dp_rfE_RAM_3__4_), .S(n684), .Y(n661) );
  MUX2NX1 U881 ( .A(dp_rfE_RAM_4__4_), .B(dp_rfE_RAM_5__4_), .S(n684), .Y(n662) );
  MUX2NX1 U882 ( .A(dp_rfE_RAM_6__4_), .B(dp_rfE_RAM_7__4_), .S(n684), .Y(n663) );
  MUX2NX1 U883 ( .A(n660), .B(n661), .S(n686), .Y(n664) );
  MUX2NX1 U884 ( .A(n662), .B(n663), .S(n686), .Y(n665) );
  MUX2NX1 U885 ( .A(dp_rfE_RAM_0__5_), .B(dp_rfE_RAM_1__5_), .S(n685), .Y(n666) );
  MUX2NX1 U886 ( .A(dp_rfE_RAM_2__5_), .B(dp_rfE_RAM_3__5_), .S(n685), .Y(n667) );
  MUX2NX1 U887 ( .A(dp_rfE_RAM_4__5_), .B(dp_rfE_RAM_5__5_), .S(n685), .Y(n668) );
  MUX2NX1 U888 ( .A(dp_rfE_RAM_6__5_), .B(dp_rfE_RAM_7__5_), .S(n685), .Y(n669) );
  MUX2NX1 U889 ( .A(n666), .B(n667), .S(n686), .Y(n670) );
  MUX2NX1 U890 ( .A(n668), .B(n669), .S(n686), .Y(n671) );
  MUX2NX1 U891 ( .A(dp_rfE_RAM_0__6_), .B(dp_rfE_RAM_1__6_), .S(n685), .Y(n672) );
  MUX2NX1 U892 ( .A(dp_rfE_RAM_2__6_), .B(dp_rfE_RAM_3__6_), .S(n685), .Y(n673) );
  MUX2NX1 U893 ( .A(dp_rfE_RAM_4__6_), .B(dp_rfE_RAM_5__6_), .S(n685), .Y(n674) );
  MUX2NX1 U894 ( .A(dp_rfE_RAM_6__6_), .B(dp_rfE_RAM_7__6_), .S(n685), .Y(n675) );
  MUX2NX1 U895 ( .A(n672), .B(n673), .S(n686), .Y(n676) );
  MUX2NX1 U896 ( .A(n674), .B(n675), .S(n686), .Y(n677) );
  MUX2NX1 U897 ( .A(dp_rfE_RAM_0__7_), .B(dp_rfE_RAM_1__7_), .S(n685), .Y(n678) );
  MUX2NX1 U898 ( .A(dp_rfE_RAM_2__7_), .B(dp_rfE_RAM_3__7_), .S(n685), .Y(n679) );
  MUX2NX1 U899 ( .A(dp_rfE_RAM_4__7_), .B(dp_rfE_RAM_5__7_), .S(n685), .Y(n680) );
  MUX2NX1 U900 ( .A(dp_rfE_RAM_6__7_), .B(dp_rfE_RAM_7__7_), .S(n685), .Y(n681) );
  MUX2NX1 U901 ( .A(n678), .B(n679), .S(n686), .Y(n682) );
  MUX2NX1 U902 ( .A(n680), .B(n681), .S(n686), .Y(n683) );
  MUX2NX1 U903 ( .A(dp_rfE_RAM_0__0_), .B(dp_rfE_RAM_1__0_), .S(n736), .Y(n687) );
  MUX2NX1 U904 ( .A(dp_rfE_RAM_2__0_), .B(dp_rfE_RAM_3__0_), .S(n736), .Y(n688) );
  MUX2NX1 U905 ( .A(dp_rfE_RAM_4__0_), .B(dp_rfE_RAM_5__0_), .S(n736), .Y(n689) );
  MUX2NX1 U906 ( .A(dp_rfE_RAM_6__0_), .B(dp_rfE_RAM_7__0_), .S(n736), .Y(n690) );
  MUX2NX1 U907 ( .A(n687), .B(n688), .S(n737), .Y(n691) );
  MUX2NX1 U908 ( .A(n689), .B(n690), .S(n737), .Y(n692) );
  MUX2NX1 U909 ( .A(dp_rfE_RAM_0__1_), .B(dp_rfE_RAM_1__1_), .S(n735), .Y(n693) );
  MUX2NX1 U910 ( .A(dp_rfE_RAM_2__1_), .B(dp_rfE_RAM_3__1_), .S(n735), .Y(n694) );
  MUX2NX1 U911 ( .A(dp_rfE_RAM_4__1_), .B(dp_rfE_RAM_5__1_), .S(n735), .Y(n695) );
  MUX2NX1 U912 ( .A(dp_rfE_RAM_6__1_), .B(dp_rfE_RAM_7__1_), .S(n735), .Y(n696) );
  MUX2NX1 U913 ( .A(n693), .B(n694), .S(n737), .Y(n697) );
  MUX2NX1 U914 ( .A(n695), .B(n696), .S(n737), .Y(n698) );
  MUX2NX1 U915 ( .A(dp_rfE_RAM_0__2_), .B(dp_rfE_RAM_1__2_), .S(n735), .Y(n699) );
  MUX2NX1 U916 ( .A(dp_rfE_RAM_2__2_), .B(dp_rfE_RAM_3__2_), .S(n735), .Y(n700) );
  MUX2NX1 U917 ( .A(dp_rfE_RAM_4__2_), .B(dp_rfE_RAM_5__2_), .S(n735), .Y(n701) );
  MUX2NX1 U918 ( .A(dp_rfE_RAM_6__2_), .B(dp_rfE_RAM_7__2_), .S(n735), .Y(n702) );
  MUX2NX1 U919 ( .A(n699), .B(n700), .S(n737), .Y(n703) );
  MUX2NX1 U920 ( .A(n701), .B(n702), .S(n737), .Y(n704) );
  MUX2NX1 U921 ( .A(dp_rfE_RAM_0__3_), .B(dp_rfE_RAM_1__3_), .S(n735), .Y(n705) );
  MUX2NX1 U922 ( .A(dp_rfE_RAM_2__3_), .B(dp_rfE_RAM_3__3_), .S(n735), .Y(n706) );
  MUX2NX1 U923 ( .A(dp_rfE_RAM_4__3_), .B(dp_rfE_RAM_5__3_), .S(n735), .Y(n707) );
  MUX2NX1 U924 ( .A(dp_rfE_RAM_6__3_), .B(dp_rfE_RAM_7__3_), .S(n735), .Y(n708) );
  MUX2NX1 U925 ( .A(n705), .B(n706), .S(n737), .Y(n709) );
  MUX2NX1 U926 ( .A(n707), .B(n708), .S(n737), .Y(n710) );
  MUX2NX1 U927 ( .A(dp_rfE_RAM_0__4_), .B(dp_rfE_RAM_1__4_), .S(n735), .Y(n711) );
  MUX2NX1 U928 ( .A(dp_rfE_RAM_2__4_), .B(dp_rfE_RAM_3__4_), .S(n735), .Y(n712) );
  MUX2NX1 U929 ( .A(dp_rfE_RAM_4__4_), .B(dp_rfE_RAM_5__4_), .S(n735), .Y(n713) );
  MUX2NX1 U930 ( .A(dp_rfE_RAM_6__4_), .B(dp_rfE_RAM_7__4_), .S(n735), .Y(n714) );
  MUX2NX1 U931 ( .A(n711), .B(n712), .S(n737), .Y(n715) );
  MUX2NX1 U932 ( .A(n713), .B(n714), .S(n737), .Y(n716) );
  MUX2NX1 U933 ( .A(dp_rfE_RAM_0__5_), .B(dp_rfE_RAM_1__5_), .S(n736), .Y(n717) );
  MUX2NX1 U934 ( .A(dp_rfE_RAM_2__5_), .B(dp_rfE_RAM_3__5_), .S(n736), .Y(n718) );
  MUX2NX1 U935 ( .A(dp_rfE_RAM_4__5_), .B(dp_rfE_RAM_5__5_), .S(n736), .Y(n719) );
  MUX2NX1 U936 ( .A(dp_rfE_RAM_6__5_), .B(dp_rfE_RAM_7__5_), .S(n736), .Y(n720) );
  MUX2NX1 U937 ( .A(n717), .B(n718), .S(n737), .Y(n721) );
  MUX2NX1 U938 ( .A(n719), .B(n720), .S(n737), .Y(n722) );
  MUX2NX1 U939 ( .A(dp_rfE_RAM_0__6_), .B(dp_rfE_RAM_1__6_), .S(n736), .Y(n723) );
  MUX2NX1 U940 ( .A(dp_rfE_RAM_2__6_), .B(dp_rfE_RAM_3__6_), .S(n736), .Y(n724) );
  MUX2NX1 U941 ( .A(dp_rfE_RAM_4__6_), .B(dp_rfE_RAM_5__6_), .S(n736), .Y(n725) );
  MUX2NX1 U942 ( .A(dp_rfE_RAM_6__6_), .B(dp_rfE_RAM_7__6_), .S(n736), .Y(n726) );
  MUX2NX1 U943 ( .A(n723), .B(n724), .S(n737), .Y(n727) );
  MUX2NX1 U944 ( .A(n725), .B(n726), .S(n737), .Y(n728) );
  MUX2NX1 U945 ( .A(dp_rfE_RAM_0__7_), .B(dp_rfE_RAM_1__7_), .S(n736), .Y(n729) );
  MUX2NX1 U946 ( .A(dp_rfE_RAM_2__7_), .B(dp_rfE_RAM_3__7_), .S(n736), .Y(n730) );
  MUX2NX1 U947 ( .A(dp_rfE_RAM_4__7_), .B(dp_rfE_RAM_5__7_), .S(n736), .Y(n731) );
  MUX2NX1 U948 ( .A(dp_rfE_RAM_6__7_), .B(dp_rfE_RAM_7__7_), .S(n736), .Y(n732) );
  MUX2NX1 U949 ( .A(n729), .B(n730), .S(n737), .Y(n733) );
  MUX2NX1 U950 ( .A(n731), .B(n732), .S(n737), .Y(n734) );
  INVX4 U951 ( .A(n745), .Y(n141) );
  INVX1 U952 ( .A(n417), .Y(n97) );
  BUFX2 U953 ( .A(dp_aluresult_0_), .Y(n738) );
  OAI21X1 U954 ( .A(n102), .B(n138), .C(n374), .Y(n739) );
  MUX2X2 U955 ( .A(n105), .B(DP_OP_50_64_8725_n71), .S(n308), .Y(
        dp_alunit_b2[2]) );
  NOR2X1 U956 ( .A(n740), .B(n742), .Y(n743) );
  NOR2X1 U957 ( .A(n743), .B(n392), .Y(n308) );
  NOR2X2 U958 ( .A(n142), .B(n745), .Y(n419) );
  NAND2X1 U959 ( .A(instr[5]), .B(n746), .Y(n747) );
  NAND2X1 U960 ( .A(n747), .B(n293), .Y(dp_nextpc[7]) );
  INVX1 U961 ( .A(instr[5]), .Y(n169) );
  NAND2X2 U962 ( .A(n286), .B(n124), .Y(n420) );
  NAND2X1 U963 ( .A(n367), .B(n368), .Y(dp_aluresult_0_) );
  INVX1 U964 ( .A(n301), .Y(n98) );
endmodule

